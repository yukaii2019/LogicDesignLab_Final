module BackGroundMemory(read_addr_color,color,clk,rst,write_en,address,w_color,block_exist,read_address,foresee,write_foresee_en,reset_foresee,store,reset_store,write_store_en);
output reg [2879:0]color;
output reg [11:0] read_addr_color;
output reg [1499:0] foresee;
output reg [299:0]store;

input clk;
input rst;
input write_en;
input [7:0]address;
input [11:0]w_color;
input [239:0]block_exist;
input [7:0]read_address;
input write_foresee_en;
input [4:0]reset_foresee;
input reset_store;
input write_store_en;

reg [2879:0]tmp_color;
reg [11:0]tmp_read_addr_color;
reg [1499:0] tmp_foresee;
reg [299:0] tmp_store;

always@(*)begin
    tmp_store = store;
    if(write_store_en)begin
        case(address)
            0 : begin tmp_store[11:0] = w_color; end
            1 : begin tmp_store[23:12] = w_color; end
            2 : begin tmp_store[35:24] = w_color; end
            3 : begin tmp_store[47:36] = w_color; end
            4 : begin tmp_store[59:48] = w_color; end
            5 : begin tmp_store[71:60] = w_color; end
            6 : begin tmp_store[83:72] = w_color; end
            7 : begin tmp_store[95:84] = w_color; end
            8 : begin tmp_store[107:96] = w_color; end
            9 : begin tmp_store[119:108] = w_color; end
            10 : begin tmp_store[131:120] = w_color; end
            11 : begin tmp_store[143:132] = w_color; end
            12 : begin tmp_store[155:144] = w_color; end
            13 : begin tmp_store[167:156] = w_color; end
            14 : begin tmp_store[179:168] = w_color; end
            15 : begin tmp_store[191:180] = w_color; end
            16 : begin tmp_store[203:192] = w_color; end
            17 : begin tmp_store[215:204] = w_color; end
            18 : begin tmp_store[227:216] = w_color; end
            19 : begin tmp_store[239:228] = w_color; end
            20 : begin tmp_store[251:240] = w_color; end
            21 : begin tmp_store[263:252] = w_color; end
            22 : begin tmp_store[275:264] = w_color; end
            23 : begin tmp_store[287:276] = w_color; end
            24 : begin tmp_store[299:288] = w_color; end
            default:begin end
        endcase
    end
    else begin
        tmp_store[11:0] = (!reset_store)?store[11:0]:12'h222;
        tmp_store[23:12] = (!reset_store)?store[23:12]:12'h111;
        tmp_store[35:24] = (!reset_store)?store[35:24]:12'h222;
        tmp_store[47:36] = (!reset_store)?store[47:36]:12'h111;
        tmp_store[59:48] = (!reset_store)?store[59:48]:12'h222;
        tmp_store[71:60] = (!reset_store)?store[71:60]:12'h111;
        tmp_store[83:72] = (!reset_store)?store[83:72]:12'h222;
        tmp_store[95:84] = (!reset_store)?store[95:84]:12'h111;
        tmp_store[107:96] = (!reset_store)?store[107:96]:12'h222;
        tmp_store[119:108] = (!reset_store)?store[119:108]:12'h111;
        tmp_store[131:120] = (!reset_store)?store[131:120]:12'h222;
        tmp_store[143:132] = (!reset_store)?store[143:132]:12'h111;
        tmp_store[155:144] = (!reset_store)?store[155:144]:12'h222;
        tmp_store[167:156] = (!reset_store)?store[167:156]:12'h111;
        tmp_store[179:168] = (!reset_store)?store[179:168]:12'h222;
        tmp_store[191:180] = (!reset_store)?store[191:180]:12'h111;
        tmp_store[203:192] = (!reset_store)?store[203:192]:12'h222;
        tmp_store[215:204] = (!reset_store)?store[215:204]:12'h111;
        tmp_store[227:216] = (!reset_store)?store[227:216]:12'h222;
        tmp_store[239:228] = (!reset_store)?store[239:228]:12'h111;
        tmp_store[251:240] = (!reset_store)?store[251:240]:12'h222;
        tmp_store[263:252] = (!reset_store)?store[263:252]:12'h111;
        tmp_store[275:264] = (!reset_store)?store[275:264]:12'h222;
        tmp_store[287:276] = (!reset_store)?store[287:276]:12'h111;
        tmp_store[299:288] = (!reset_store)?store[299:288]:12'h222;
    end
end
always@(*)begin
    tmp_foresee = foresee;
    if(write_foresee_en)begin
        case(address)
            0 : begin tmp_foresee[11:0] = w_color; end
            1 : begin tmp_foresee[23:12] = w_color; end
            2 : begin tmp_foresee[35:24] = w_color; end
            3 : begin tmp_foresee[47:36] = w_color; end
            4 : begin tmp_foresee[59:48] = w_color; end
            5 : begin tmp_foresee[71:60] = w_color; end
            6 : begin tmp_foresee[83:72] = w_color; end
            7 : begin tmp_foresee[95:84] = w_color; end
            8 : begin tmp_foresee[107:96] = w_color; end
            9 : begin tmp_foresee[119:108] = w_color; end
            10 : begin tmp_foresee[131:120] = w_color; end
            11 : begin tmp_foresee[143:132] = w_color; end
            12 : begin tmp_foresee[155:144] = w_color; end
            13 : begin tmp_foresee[167:156] = w_color; end
            14 : begin tmp_foresee[179:168] = w_color; end
            15 : begin tmp_foresee[191:180] = w_color; end
            16 : begin tmp_foresee[203:192] = w_color; end
            17 : begin tmp_foresee[215:204] = w_color; end
            18 : begin tmp_foresee[227:216] = w_color; end
            19 : begin tmp_foresee[239:228] = w_color; end
            20 : begin tmp_foresee[251:240] = w_color; end
            21 : begin tmp_foresee[263:252] = w_color; end
            22 : begin tmp_foresee[275:264] = w_color; end
            23 : begin tmp_foresee[287:276] = w_color; end
            24 : begin tmp_foresee[299:288] = w_color; end
            25 : begin tmp_foresee[311:300] = w_color; end
            26 : begin tmp_foresee[323:312] = w_color; end
            27 : begin tmp_foresee[335:324] = w_color; end
            28 : begin tmp_foresee[347:336] = w_color; end
            29 : begin tmp_foresee[359:348] = w_color; end
            30 : begin tmp_foresee[371:360] = w_color; end
            31 : begin tmp_foresee[383:372] = w_color; end
            32 : begin tmp_foresee[395:384] = w_color; end
            33 : begin tmp_foresee[407:396] = w_color; end
            34 : begin tmp_foresee[419:408] = w_color; end
            35 : begin tmp_foresee[431:420] = w_color; end
            36 : begin tmp_foresee[443:432] = w_color; end
            37 : begin tmp_foresee[455:444] = w_color; end
            38 : begin tmp_foresee[467:456] = w_color; end
            39 : begin tmp_foresee[479:468] = w_color; end
            40 : begin tmp_foresee[491:480] = w_color; end
            41 : begin tmp_foresee[503:492] = w_color; end
            42 : begin tmp_foresee[515:504] = w_color; end
            43 : begin tmp_foresee[527:516] = w_color; end
            44 : begin tmp_foresee[539:528] = w_color; end
            45 : begin tmp_foresee[551:540] = w_color; end
            46 : begin tmp_foresee[563:552] = w_color; end
            47 : begin tmp_foresee[575:564] = w_color; end
            48 : begin tmp_foresee[587:576] = w_color; end
            49 : begin tmp_foresee[599:588] = w_color; end
            50 : begin tmp_foresee[611:600] = w_color; end
            51 : begin tmp_foresee[623:612] = w_color; end
            52 : begin tmp_foresee[635:624] = w_color; end
            53 : begin tmp_foresee[647:636] = w_color; end
            54 : begin tmp_foresee[659:648] = w_color; end
            55 : begin tmp_foresee[671:660] = w_color; end
            56 : begin tmp_foresee[683:672] = w_color; end
            57 : begin tmp_foresee[695:684] = w_color; end
            58 : begin tmp_foresee[707:696] = w_color; end
            59 : begin tmp_foresee[719:708] = w_color; end
            60 : begin tmp_foresee[731:720] = w_color; end
            61 : begin tmp_foresee[743:732] = w_color; end
            62 : begin tmp_foresee[755:744] = w_color; end
            63 : begin tmp_foresee[767:756] = w_color; end
            64 : begin tmp_foresee[779:768] = w_color; end
            65 : begin tmp_foresee[791:780] = w_color; end
            66 : begin tmp_foresee[803:792] = w_color; end
            67 : begin tmp_foresee[815:804] = w_color; end
            68 : begin tmp_foresee[827:816] = w_color; end
            69 : begin tmp_foresee[839:828] = w_color; end
            70 : begin tmp_foresee[851:840] = w_color; end
            71 : begin tmp_foresee[863:852] = w_color; end
            72 : begin tmp_foresee[875:864] = w_color; end
            73 : begin tmp_foresee[887:876] = w_color; end
            74 : begin tmp_foresee[899:888] = w_color; end
            75 : begin tmp_foresee[911:900] = w_color; end
            76 : begin tmp_foresee[923:912] = w_color; end
            77 : begin tmp_foresee[935:924] = w_color; end
            78 : begin tmp_foresee[947:936] = w_color; end
            79 : begin tmp_foresee[959:948] = w_color; end
            80 : begin tmp_foresee[971:960] = w_color; end
            81 : begin tmp_foresee[983:972] = w_color; end
            82 : begin tmp_foresee[995:984] = w_color; end
            83 : begin tmp_foresee[1007:996] = w_color; end
            84 : begin tmp_foresee[1019:1008] = w_color; end
            85 : begin tmp_foresee[1031:1020] = w_color; end
            86 : begin tmp_foresee[1043:1032] = w_color; end
            87 : begin tmp_foresee[1055:1044] = w_color; end
            88 : begin tmp_foresee[1067:1056] = w_color; end
            89 : begin tmp_foresee[1079:1068] = w_color; end
            90 : begin tmp_foresee[1091:1080] = w_color; end
            91 : begin tmp_foresee[1103:1092] = w_color; end
            92 : begin tmp_foresee[1115:1104] = w_color; end
            93 : begin tmp_foresee[1127:1116] = w_color; end
            94 : begin tmp_foresee[1139:1128] = w_color; end
            95 : begin tmp_foresee[1151:1140] = w_color; end
            96 : begin tmp_foresee[1163:1152] = w_color; end
            97 : begin tmp_foresee[1175:1164] = w_color; end
            98 : begin tmp_foresee[1187:1176] = w_color; end
            99 : begin tmp_foresee[1199:1188] = w_color; end
            100 : begin tmp_foresee[1211:1200] = w_color; end
            101 : begin tmp_foresee[1223:1212] = w_color; end
            102 : begin tmp_foresee[1235:1224] = w_color; end
            103 : begin tmp_foresee[1247:1236] = w_color; end
            104 : begin tmp_foresee[1259:1248] = w_color; end
            105 : begin tmp_foresee[1271:1260] = w_color; end
            106 : begin tmp_foresee[1283:1272] = w_color; end
            107 : begin tmp_foresee[1295:1284] = w_color; end
            108 : begin tmp_foresee[1307:1296] = w_color; end
            109 : begin tmp_foresee[1319:1308] = w_color; end
            110 : begin tmp_foresee[1331:1320] = w_color; end
            111 : begin tmp_foresee[1343:1332] = w_color; end
            112 : begin tmp_foresee[1355:1344] = w_color; end
            113 : begin tmp_foresee[1367:1356] = w_color; end
            114 : begin tmp_foresee[1379:1368] = w_color; end
            115 : begin tmp_foresee[1391:1380] = w_color; end
            116 : begin tmp_foresee[1403:1392] = w_color; end
            117 : begin tmp_foresee[1415:1404] = w_color; end
            118 : begin tmp_foresee[1427:1416] = w_color; end
            119 : begin tmp_foresee[1439:1428] = w_color; end
            120 : begin tmp_foresee[1451:1440] = w_color; end
            121 : begin tmp_foresee[1463:1452] = w_color; end
            122 : begin tmp_foresee[1475:1464] = w_color; end
            123 : begin tmp_foresee[1487:1476] = w_color; end
            124 : begin tmp_foresee[1499:1488] = w_color; end
            default:begin end
        endcase
    end
    else begin
tmp_foresee[11:0] = (!reset_foresee[0])?foresee[11:0]:12'h222;
tmp_foresee[23:12] = (!reset_foresee[0])?foresee[23:12]:12'h111;
tmp_foresee[35:24] = (!reset_foresee[0])?foresee[35:24]:12'h222;
tmp_foresee[47:36] = (!reset_foresee[0])?foresee[47:36]:12'h111;
tmp_foresee[59:48] = (!reset_foresee[0])?foresee[59:48]:12'h222;
tmp_foresee[71:60] = (!reset_foresee[0])?foresee[71:60]:12'h111;
tmp_foresee[83:72] = (!reset_foresee[0])?foresee[83:72]:12'h222;
tmp_foresee[95:84] = (!reset_foresee[0])?foresee[95:84]:12'h111;
tmp_foresee[107:96] = (!reset_foresee[0])?foresee[107:96]:12'h222;
tmp_foresee[119:108] = (!reset_foresee[0])?foresee[119:108]:12'h111;
tmp_foresee[131:120] = (!reset_foresee[0])?foresee[131:120]:12'h222;
tmp_foresee[143:132] = (!reset_foresee[0])?foresee[143:132]:12'h111;
tmp_foresee[155:144] = (!reset_foresee[0])?foresee[155:144]:12'h222;
tmp_foresee[167:156] = (!reset_foresee[0])?foresee[167:156]:12'h111;
tmp_foresee[179:168] = (!reset_foresee[0])?foresee[179:168]:12'h222;
tmp_foresee[191:180] = (!reset_foresee[0])?foresee[191:180]:12'h111;
tmp_foresee[203:192] = (!reset_foresee[0])?foresee[203:192]:12'h222;
tmp_foresee[215:204] = (!reset_foresee[0])?foresee[215:204]:12'h111;
tmp_foresee[227:216] = (!reset_foresee[0])?foresee[227:216]:12'h222;
tmp_foresee[239:228] = (!reset_foresee[0])?foresee[239:228]:12'h111;
tmp_foresee[251:240] = (!reset_foresee[0])?foresee[251:240]:12'h222;
tmp_foresee[263:252] = (!reset_foresee[0])?foresee[263:252]:12'h111;
tmp_foresee[275:264] = (!reset_foresee[0])?foresee[275:264]:12'h222;
tmp_foresee[287:276] = (!reset_foresee[0])?foresee[287:276]:12'h111;
tmp_foresee[299:288] = (!reset_foresee[0])?foresee[299:288]:12'h222;
tmp_foresee[311:300] = (!reset_foresee[1])?foresee[311:300]:12'h111;
tmp_foresee[323:312] = (!reset_foresee[1])?foresee[323:312]:12'h222;
tmp_foresee[335:324] = (!reset_foresee[1])?foresee[335:324]:12'h111;
tmp_foresee[347:336] = (!reset_foresee[1])?foresee[347:336]:12'h222;
tmp_foresee[359:348] = (!reset_foresee[1])?foresee[359:348]:12'h111;
tmp_foresee[371:360] = (!reset_foresee[1])?foresee[371:360]:12'h222;
tmp_foresee[383:372] = (!reset_foresee[1])?foresee[383:372]:12'h111;
tmp_foresee[395:384] = (!reset_foresee[1])?foresee[395:384]:12'h222;
tmp_foresee[407:396] = (!reset_foresee[1])?foresee[407:396]:12'h111;
tmp_foresee[419:408] = (!reset_foresee[1])?foresee[419:408]:12'h222;
tmp_foresee[431:420] = (!reset_foresee[1])?foresee[431:420]:12'h111;
tmp_foresee[443:432] = (!reset_foresee[1])?foresee[443:432]:12'h222;
tmp_foresee[455:444] = (!reset_foresee[1])?foresee[455:444]:12'h111;
tmp_foresee[467:456] = (!reset_foresee[1])?foresee[467:456]:12'h222;
tmp_foresee[479:468] = (!reset_foresee[1])?foresee[479:468]:12'h111;
tmp_foresee[491:480] = (!reset_foresee[1])?foresee[491:480]:12'h222;
tmp_foresee[503:492] = (!reset_foresee[1])?foresee[503:492]:12'h111;
tmp_foresee[515:504] = (!reset_foresee[1])?foresee[515:504]:12'h222;
tmp_foresee[527:516] = (!reset_foresee[1])?foresee[527:516]:12'h111;
tmp_foresee[539:528] = (!reset_foresee[1])?foresee[539:528]:12'h222;
tmp_foresee[551:540] = (!reset_foresee[1])?foresee[551:540]:12'h111;
tmp_foresee[563:552] = (!reset_foresee[1])?foresee[563:552]:12'h222;
tmp_foresee[575:564] = (!reset_foresee[1])?foresee[575:564]:12'h111;
tmp_foresee[587:576] = (!reset_foresee[1])?foresee[587:576]:12'h222;
tmp_foresee[599:588] = (!reset_foresee[1])?foresee[599:588]:12'h111;
tmp_foresee[611:600] = (!reset_foresee[2])?foresee[611:600]:12'h222;
tmp_foresee[623:612] = (!reset_foresee[2])?foresee[623:612]:12'h111;
tmp_foresee[635:624] = (!reset_foresee[2])?foresee[635:624]:12'h222;
tmp_foresee[647:636] = (!reset_foresee[2])?foresee[647:636]:12'h111;
tmp_foresee[659:648] = (!reset_foresee[2])?foresee[659:648]:12'h222;
tmp_foresee[671:660] = (!reset_foresee[2])?foresee[671:660]:12'h111;
tmp_foresee[683:672] = (!reset_foresee[2])?foresee[683:672]:12'h222;
tmp_foresee[695:684] = (!reset_foresee[2])?foresee[695:684]:12'h111;
tmp_foresee[707:696] = (!reset_foresee[2])?foresee[707:696]:12'h222;
tmp_foresee[719:708] = (!reset_foresee[2])?foresee[719:708]:12'h111;
tmp_foresee[731:720] = (!reset_foresee[2])?foresee[731:720]:12'h222;
tmp_foresee[743:732] = (!reset_foresee[2])?foresee[743:732]:12'h111;
tmp_foresee[755:744] = (!reset_foresee[2])?foresee[755:744]:12'h222;
tmp_foresee[767:756] = (!reset_foresee[2])?foresee[767:756]:12'h111;
tmp_foresee[779:768] = (!reset_foresee[2])?foresee[779:768]:12'h222;
tmp_foresee[791:780] = (!reset_foresee[2])?foresee[791:780]:12'h111;
tmp_foresee[803:792] = (!reset_foresee[2])?foresee[803:792]:12'h222;
tmp_foresee[815:804] = (!reset_foresee[2])?foresee[815:804]:12'h111;
tmp_foresee[827:816] = (!reset_foresee[2])?foresee[827:816]:12'h222;
tmp_foresee[839:828] = (!reset_foresee[2])?foresee[839:828]:12'h111;
tmp_foresee[851:840] = (!reset_foresee[2])?foresee[851:840]:12'h222;
tmp_foresee[863:852] = (!reset_foresee[2])?foresee[863:852]:12'h111;
tmp_foresee[875:864] = (!reset_foresee[2])?foresee[875:864]:12'h222;
tmp_foresee[887:876] = (!reset_foresee[2])?foresee[887:876]:12'h111;
tmp_foresee[899:888] = (!reset_foresee[2])?foresee[899:888]:12'h222;
tmp_foresee[911:900] = (!reset_foresee[3])?foresee[911:900]:12'h111;
tmp_foresee[923:912] = (!reset_foresee[3])?foresee[923:912]:12'h222;
tmp_foresee[935:924] = (!reset_foresee[3])?foresee[935:924]:12'h111;
tmp_foresee[947:936] = (!reset_foresee[3])?foresee[947:936]:12'h222;
tmp_foresee[959:948] = (!reset_foresee[3])?foresee[959:948]:12'h111;
tmp_foresee[971:960] = (!reset_foresee[3])?foresee[971:960]:12'h222;
tmp_foresee[983:972] = (!reset_foresee[3])?foresee[983:972]:12'h111;
tmp_foresee[995:984] = (!reset_foresee[3])?foresee[995:984]:12'h222;
tmp_foresee[1007:996] = (!reset_foresee[3])?foresee[1007:996]:12'h111;
tmp_foresee[1019:1008] = (!reset_foresee[3])?foresee[1019:1008]:12'h222;
tmp_foresee[1031:1020] = (!reset_foresee[3])?foresee[1031:1020]:12'h111;
tmp_foresee[1043:1032] = (!reset_foresee[3])?foresee[1043:1032]:12'h222;
tmp_foresee[1055:1044] = (!reset_foresee[3])?foresee[1055:1044]:12'h111;
tmp_foresee[1067:1056] = (!reset_foresee[3])?foresee[1067:1056]:12'h222;
tmp_foresee[1079:1068] = (!reset_foresee[3])?foresee[1079:1068]:12'h111;
tmp_foresee[1091:1080] = (!reset_foresee[3])?foresee[1091:1080]:12'h222;
tmp_foresee[1103:1092] = (!reset_foresee[3])?foresee[1103:1092]:12'h111;
tmp_foresee[1115:1104] = (!reset_foresee[3])?foresee[1115:1104]:12'h222;
tmp_foresee[1127:1116] = (!reset_foresee[3])?foresee[1127:1116]:12'h111;
tmp_foresee[1139:1128] = (!reset_foresee[3])?foresee[1139:1128]:12'h222;
tmp_foresee[1151:1140] = (!reset_foresee[3])?foresee[1151:1140]:12'h111;
tmp_foresee[1163:1152] = (!reset_foresee[3])?foresee[1163:1152]:12'h222;
tmp_foresee[1175:1164] = (!reset_foresee[3])?foresee[1175:1164]:12'h111;
tmp_foresee[1187:1176] = (!reset_foresee[3])?foresee[1187:1176]:12'h222;
tmp_foresee[1199:1188] = (!reset_foresee[3])?foresee[1199:1188]:12'h111;
tmp_foresee[1211:1200] = (!reset_foresee[4])?foresee[1211:1200]:12'h222;
tmp_foresee[1223:1212] = (!reset_foresee[4])?foresee[1223:1212]:12'h111;
tmp_foresee[1235:1224] = (!reset_foresee[4])?foresee[1235:1224]:12'h222;
tmp_foresee[1247:1236] = (!reset_foresee[4])?foresee[1247:1236]:12'h111;
tmp_foresee[1259:1248] = (!reset_foresee[4])?foresee[1259:1248]:12'h222;
tmp_foresee[1271:1260] = (!reset_foresee[4])?foresee[1271:1260]:12'h111;
tmp_foresee[1283:1272] = (!reset_foresee[4])?foresee[1283:1272]:12'h222;
tmp_foresee[1295:1284] = (!reset_foresee[4])?foresee[1295:1284]:12'h111;
tmp_foresee[1307:1296] = (!reset_foresee[4])?foresee[1307:1296]:12'h222;
tmp_foresee[1319:1308] = (!reset_foresee[4])?foresee[1319:1308]:12'h111;
tmp_foresee[1331:1320] = (!reset_foresee[4])?foresee[1331:1320]:12'h222;
tmp_foresee[1343:1332] = (!reset_foresee[4])?foresee[1343:1332]:12'h111;
tmp_foresee[1355:1344] = (!reset_foresee[4])?foresee[1355:1344]:12'h222;
tmp_foresee[1367:1356] = (!reset_foresee[4])?foresee[1367:1356]:12'h111;
tmp_foresee[1379:1368] = (!reset_foresee[4])?foresee[1379:1368]:12'h222;
tmp_foresee[1391:1380] = (!reset_foresee[4])?foresee[1391:1380]:12'h111;
tmp_foresee[1403:1392] = (!reset_foresee[4])?foresee[1403:1392]:12'h222;
tmp_foresee[1415:1404] = (!reset_foresee[4])?foresee[1415:1404]:12'h111;
tmp_foresee[1427:1416] = (!reset_foresee[4])?foresee[1427:1416]:12'h222;
tmp_foresee[1439:1428] = (!reset_foresee[4])?foresee[1439:1428]:12'h111;
tmp_foresee[1451:1440] = (!reset_foresee[4])?foresee[1451:1440]:12'h222;
tmp_foresee[1463:1452] = (!reset_foresee[4])?foresee[1463:1452]:12'h111;
tmp_foresee[1475:1464] = (!reset_foresee[4])?foresee[1475:1464]:12'h222;
tmp_foresee[1487:1476] = (!reset_foresee[4])?foresee[1487:1476]:12'h111;
tmp_foresee[1499:1488] = (!reset_foresee[4])?foresee[1499:1488]:12'h222;

    end
end
always@(*)begin
    tmp_read_addr_color = read_addr_color;
    case(read_address)
        0 : begin tmp_read_addr_color = color[11:0]; end
        1 : begin tmp_read_addr_color = color[23:12]; end
        2 : begin tmp_read_addr_color = color[35:24]; end
        3 : begin tmp_read_addr_color = color[47:36]; end
        4 : begin tmp_read_addr_color = color[59:48]; end
        5 : begin tmp_read_addr_color = color[71:60]; end
        6 : begin tmp_read_addr_color = color[83:72]; end
        7 : begin tmp_read_addr_color = color[95:84]; end
        8 : begin tmp_read_addr_color = color[107:96]; end
        9 : begin tmp_read_addr_color = color[119:108]; end
        10 : begin tmp_read_addr_color = color[131:120]; end
        11 : begin tmp_read_addr_color = color[143:132]; end
        12 : begin tmp_read_addr_color = color[155:144]; end
        13 : begin tmp_read_addr_color = color[167:156]; end
        14 : begin tmp_read_addr_color = color[179:168]; end
        15 : begin tmp_read_addr_color = color[191:180]; end
        16 : begin tmp_read_addr_color = color[203:192]; end
        17 : begin tmp_read_addr_color = color[215:204]; end
        18 : begin tmp_read_addr_color = color[227:216]; end
        19 : begin tmp_read_addr_color = color[239:228]; end
        20 : begin tmp_read_addr_color = color[251:240]; end
        21 : begin tmp_read_addr_color = color[263:252]; end
        22 : begin tmp_read_addr_color = color[275:264]; end
        23 : begin tmp_read_addr_color = color[287:276]; end
        24 : begin tmp_read_addr_color = color[299:288]; end
        25 : begin tmp_read_addr_color = color[311:300]; end
        26 : begin tmp_read_addr_color = color[323:312]; end
        27 : begin tmp_read_addr_color = color[335:324]; end
        28 : begin tmp_read_addr_color = color[347:336]; end
        29 : begin tmp_read_addr_color = color[359:348]; end
        30 : begin tmp_read_addr_color = color[371:360]; end
        31 : begin tmp_read_addr_color = color[383:372]; end
        32 : begin tmp_read_addr_color = color[395:384]; end
        33 : begin tmp_read_addr_color = color[407:396]; end
        34 : begin tmp_read_addr_color = color[419:408]; end
        35 : begin tmp_read_addr_color = color[431:420]; end
        36 : begin tmp_read_addr_color = color[443:432]; end
        37 : begin tmp_read_addr_color = color[455:444]; end
        38 : begin tmp_read_addr_color = color[467:456]; end
        39 : begin tmp_read_addr_color = color[479:468]; end
        40 : begin tmp_read_addr_color = color[491:480]; end
        41 : begin tmp_read_addr_color = color[503:492]; end
        42 : begin tmp_read_addr_color = color[515:504]; end
        43 : begin tmp_read_addr_color = color[527:516]; end
        44 : begin tmp_read_addr_color = color[539:528]; end
        45 : begin tmp_read_addr_color = color[551:540]; end
        46 : begin tmp_read_addr_color = color[563:552]; end
        47 : begin tmp_read_addr_color = color[575:564]; end
        48 : begin tmp_read_addr_color = color[587:576]; end
        49 : begin tmp_read_addr_color = color[599:588]; end
        50 : begin tmp_read_addr_color = color[611:600]; end
        51 : begin tmp_read_addr_color = color[623:612]; end
        52 : begin tmp_read_addr_color = color[635:624]; end
        53 : begin tmp_read_addr_color = color[647:636]; end
        54 : begin tmp_read_addr_color = color[659:648]; end
        55 : begin tmp_read_addr_color = color[671:660]; end
        56 : begin tmp_read_addr_color = color[683:672]; end
        57 : begin tmp_read_addr_color = color[695:684]; end
        58 : begin tmp_read_addr_color = color[707:696]; end
        59 : begin tmp_read_addr_color = color[719:708]; end
        60 : begin tmp_read_addr_color = color[731:720]; end
        61 : begin tmp_read_addr_color = color[743:732]; end
        62 : begin tmp_read_addr_color = color[755:744]; end
        63 : begin tmp_read_addr_color = color[767:756]; end
        64 : begin tmp_read_addr_color = color[779:768]; end
        65 : begin tmp_read_addr_color = color[791:780]; end
        66 : begin tmp_read_addr_color = color[803:792]; end
        67 : begin tmp_read_addr_color = color[815:804]; end
        68 : begin tmp_read_addr_color = color[827:816]; end
        69 : begin tmp_read_addr_color = color[839:828]; end
        70 : begin tmp_read_addr_color = color[851:840]; end
        71 : begin tmp_read_addr_color = color[863:852]; end
        72 : begin tmp_read_addr_color = color[875:864]; end
        73 : begin tmp_read_addr_color = color[887:876]; end
        74 : begin tmp_read_addr_color = color[899:888]; end
        75 : begin tmp_read_addr_color = color[911:900]; end
        76 : begin tmp_read_addr_color = color[923:912]; end
        77 : begin tmp_read_addr_color = color[935:924]; end
        78 : begin tmp_read_addr_color = color[947:936]; end
        79 : begin tmp_read_addr_color = color[959:948]; end
        80 : begin tmp_read_addr_color = color[971:960]; end
        81 : begin tmp_read_addr_color = color[983:972]; end
        82 : begin tmp_read_addr_color = color[995:984]; end
        83 : begin tmp_read_addr_color = color[1007:996]; end
        84 : begin tmp_read_addr_color = color[1019:1008]; end
        85 : begin tmp_read_addr_color = color[1031:1020]; end
        86 : begin tmp_read_addr_color = color[1043:1032]; end
        87 : begin tmp_read_addr_color = color[1055:1044]; end
        88 : begin tmp_read_addr_color = color[1067:1056]; end
        89 : begin tmp_read_addr_color = color[1079:1068]; end
        90 : begin tmp_read_addr_color = color[1091:1080]; end
        91 : begin tmp_read_addr_color = color[1103:1092]; end
        92 : begin tmp_read_addr_color = color[1115:1104]; end
        93 : begin tmp_read_addr_color = color[1127:1116]; end
        94 : begin tmp_read_addr_color = color[1139:1128]; end
        95 : begin tmp_read_addr_color = color[1151:1140]; end
        96 : begin tmp_read_addr_color = color[1163:1152]; end
        97 : begin tmp_read_addr_color = color[1175:1164]; end
        98 : begin tmp_read_addr_color = color[1187:1176]; end
        99 : begin tmp_read_addr_color = color[1199:1188]; end
        100 : begin tmp_read_addr_color = color[1211:1200]; end
        101 : begin tmp_read_addr_color = color[1223:1212]; end
        102 : begin tmp_read_addr_color = color[1235:1224]; end
        103 : begin tmp_read_addr_color = color[1247:1236]; end
        104 : begin tmp_read_addr_color = color[1259:1248]; end
        105 : begin tmp_read_addr_color = color[1271:1260]; end
        106 : begin tmp_read_addr_color = color[1283:1272]; end
        107 : begin tmp_read_addr_color = color[1295:1284]; end
        108 : begin tmp_read_addr_color = color[1307:1296]; end
        109 : begin tmp_read_addr_color = color[1319:1308]; end
        110 : begin tmp_read_addr_color = color[1331:1320]; end
        111 : begin tmp_read_addr_color = color[1343:1332]; end
        112 : begin tmp_read_addr_color = color[1355:1344]; end
        113 : begin tmp_read_addr_color = color[1367:1356]; end
        114 : begin tmp_read_addr_color = color[1379:1368]; end
        115 : begin tmp_read_addr_color = color[1391:1380]; end
        116 : begin tmp_read_addr_color = color[1403:1392]; end
        117 : begin tmp_read_addr_color = color[1415:1404]; end
        118 : begin tmp_read_addr_color = color[1427:1416]; end
        119 : begin tmp_read_addr_color = color[1439:1428]; end
        120 : begin tmp_read_addr_color = color[1451:1440]; end
        121 : begin tmp_read_addr_color = color[1463:1452]; end
        122 : begin tmp_read_addr_color = color[1475:1464]; end
        123 : begin tmp_read_addr_color = color[1487:1476]; end
        124 : begin tmp_read_addr_color = color[1499:1488]; end
        125 : begin tmp_read_addr_color = color[1511:1500]; end
        126 : begin tmp_read_addr_color = color[1523:1512]; end
        127 : begin tmp_read_addr_color = color[1535:1524]; end
        128 : begin tmp_read_addr_color = color[1547:1536]; end
        129 : begin tmp_read_addr_color = color[1559:1548]; end
        130 : begin tmp_read_addr_color = color[1571:1560]; end
        131 : begin tmp_read_addr_color = color[1583:1572]; end
        132 : begin tmp_read_addr_color = color[1595:1584]; end
        133 : begin tmp_read_addr_color = color[1607:1596]; end
        134 : begin tmp_read_addr_color = color[1619:1608]; end
        135 : begin tmp_read_addr_color = color[1631:1620]; end
        136 : begin tmp_read_addr_color = color[1643:1632]; end
        137 : begin tmp_read_addr_color = color[1655:1644]; end
        138 : begin tmp_read_addr_color = color[1667:1656]; end
        139 : begin tmp_read_addr_color = color[1679:1668]; end
        140 : begin tmp_read_addr_color = color[1691:1680]; end
        141 : begin tmp_read_addr_color = color[1703:1692]; end
        142 : begin tmp_read_addr_color = color[1715:1704]; end
        143 : begin tmp_read_addr_color = color[1727:1716]; end
        144 : begin tmp_read_addr_color = color[1739:1728]; end
        145 : begin tmp_read_addr_color = color[1751:1740]; end
        146 : begin tmp_read_addr_color = color[1763:1752]; end
        147 : begin tmp_read_addr_color = color[1775:1764]; end
        148 : begin tmp_read_addr_color = color[1787:1776]; end
        149 : begin tmp_read_addr_color = color[1799:1788]; end
        150 : begin tmp_read_addr_color = color[1811:1800]; end
        151 : begin tmp_read_addr_color = color[1823:1812]; end
        152 : begin tmp_read_addr_color = color[1835:1824]; end
        153 : begin tmp_read_addr_color = color[1847:1836]; end
        154 : begin tmp_read_addr_color = color[1859:1848]; end
        155 : begin tmp_read_addr_color = color[1871:1860]; end
        156 : begin tmp_read_addr_color = color[1883:1872]; end
        157 : begin tmp_read_addr_color = color[1895:1884]; end
        158 : begin tmp_read_addr_color = color[1907:1896]; end
        159 : begin tmp_read_addr_color = color[1919:1908]; end
        160 : begin tmp_read_addr_color = color[1931:1920]; end
        161 : begin tmp_read_addr_color = color[1943:1932]; end
        162 : begin tmp_read_addr_color = color[1955:1944]; end
        163 : begin tmp_read_addr_color = color[1967:1956]; end
        164 : begin tmp_read_addr_color = color[1979:1968]; end
        165 : begin tmp_read_addr_color = color[1991:1980]; end
        166 : begin tmp_read_addr_color = color[2003:1992]; end
        167 : begin tmp_read_addr_color = color[2015:2004]; end
        168 : begin tmp_read_addr_color = color[2027:2016]; end
        169 : begin tmp_read_addr_color = color[2039:2028]; end
        170 : begin tmp_read_addr_color = color[2051:2040]; end
        171 : begin tmp_read_addr_color = color[2063:2052]; end
        172 : begin tmp_read_addr_color = color[2075:2064]; end
        173 : begin tmp_read_addr_color = color[2087:2076]; end
        174 : begin tmp_read_addr_color = color[2099:2088]; end
        175 : begin tmp_read_addr_color = color[2111:2100]; end
        176 : begin tmp_read_addr_color = color[2123:2112]; end
        177 : begin tmp_read_addr_color = color[2135:2124]; end
        178 : begin tmp_read_addr_color = color[2147:2136]; end
        179 : begin tmp_read_addr_color = color[2159:2148]; end
        180 : begin tmp_read_addr_color = color[2171:2160]; end
        181 : begin tmp_read_addr_color = color[2183:2172]; end
        182 : begin tmp_read_addr_color = color[2195:2184]; end
        183 : begin tmp_read_addr_color = color[2207:2196]; end
        184 : begin tmp_read_addr_color = color[2219:2208]; end
        185 : begin tmp_read_addr_color = color[2231:2220]; end
        186 : begin tmp_read_addr_color = color[2243:2232]; end
        187 : begin tmp_read_addr_color = color[2255:2244]; end
        188 : begin tmp_read_addr_color = color[2267:2256]; end
        189 : begin tmp_read_addr_color = color[2279:2268]; end
        190 : begin tmp_read_addr_color = color[2291:2280]; end
        191 : begin tmp_read_addr_color = color[2303:2292]; end
        192 : begin tmp_read_addr_color = color[2315:2304]; end
        193 : begin tmp_read_addr_color = color[2327:2316]; end
        194 : begin tmp_read_addr_color = color[2339:2328]; end
        195 : begin tmp_read_addr_color = color[2351:2340]; end
        196 : begin tmp_read_addr_color = color[2363:2352]; end
        197 : begin tmp_read_addr_color = color[2375:2364]; end
        198 : begin tmp_read_addr_color = color[2387:2376]; end
        199 : begin tmp_read_addr_color = color[2399:2388]; end
        200 : begin tmp_read_addr_color = color[2411:2400]; end
        201 : begin tmp_read_addr_color = color[2423:2412]; end
        202 : begin tmp_read_addr_color = color[2435:2424]; end
        203 : begin tmp_read_addr_color = color[2447:2436]; end
        204 : begin tmp_read_addr_color = color[2459:2448]; end
        205 : begin tmp_read_addr_color = color[2471:2460]; end
        206 : begin tmp_read_addr_color = color[2483:2472]; end
        207 : begin tmp_read_addr_color = color[2495:2484]; end
        208 : begin tmp_read_addr_color = color[2507:2496]; end
        209 : begin tmp_read_addr_color = color[2519:2508]; end
        210 : begin tmp_read_addr_color = color[2531:2520]; end
        211 : begin tmp_read_addr_color = color[2543:2532]; end
        212 : begin tmp_read_addr_color = color[2555:2544]; end
        213 : begin tmp_read_addr_color = color[2567:2556]; end
        214 : begin tmp_read_addr_color = color[2579:2568]; end
        215 : begin tmp_read_addr_color = color[2591:2580]; end
        216 : begin tmp_read_addr_color = color[2603:2592]; end
        217 : begin tmp_read_addr_color = color[2615:2604]; end
        218 : begin tmp_read_addr_color = color[2627:2616]; end
        219 : begin tmp_read_addr_color = color[2639:2628]; end
        220 : begin tmp_read_addr_color = color[2651:2640]; end
        221 : begin tmp_read_addr_color = color[2663:2652]; end
        222 : begin tmp_read_addr_color = color[2675:2664]; end
        223 : begin tmp_read_addr_color = color[2687:2676]; end
        224 : begin tmp_read_addr_color = color[2699:2688]; end
        225 : begin tmp_read_addr_color = color[2711:2700]; end
        226 : begin tmp_read_addr_color = color[2723:2712]; end
        227 : begin tmp_read_addr_color = color[2735:2724]; end
        228 : begin tmp_read_addr_color = color[2747:2736]; end
        229 : begin tmp_read_addr_color = color[2759:2748]; end
        230 : begin tmp_read_addr_color = color[2771:2760]; end
        231 : begin tmp_read_addr_color = color[2783:2772]; end
        232 : begin tmp_read_addr_color = color[2795:2784]; end
        233 : begin tmp_read_addr_color = color[2807:2796]; end
        234 : begin tmp_read_addr_color = color[2819:2808]; end
        235 : begin tmp_read_addr_color = color[2831:2820]; end
        236 : begin tmp_read_addr_color = color[2843:2832]; end
        237 : begin tmp_read_addr_color = color[2855:2844]; end
        238 : begin tmp_read_addr_color = color[2867:2856]; end
        239 : begin tmp_read_addr_color = color[2879:2868]; end
    endcase
end
always@(*)begin
    tmp_color = color;
    if(write_en)begin
        case(address)
            0 : begin tmp_color[11:0] = w_color; end
            1 : begin tmp_color[23:12] = w_color; end
            2 : begin tmp_color[35:24] = w_color; end
            3 : begin tmp_color[47:36] = w_color; end
            4 : begin tmp_color[59:48] = w_color; end
            5 : begin tmp_color[71:60] = w_color; end
            6 : begin tmp_color[83:72] = w_color; end
            7 : begin tmp_color[95:84] = w_color; end
            8 : begin tmp_color[107:96] = w_color; end
            9 : begin tmp_color[119:108] = w_color; end
            10 : begin tmp_color[131:120] = w_color; end
            11 : begin tmp_color[143:132] = w_color; end
            12 : begin tmp_color[155:144] = w_color; end
            13 : begin tmp_color[167:156] = w_color; end
            14 : begin tmp_color[179:168] = w_color; end
            15 : begin tmp_color[191:180] = w_color; end
            16 : begin tmp_color[203:192] = w_color; end
            17 : begin tmp_color[215:204] = w_color; end
            18 : begin tmp_color[227:216] = w_color; end
            19 : begin tmp_color[239:228] = w_color; end
            20 : begin tmp_color[251:240] = w_color; end
            21 : begin tmp_color[263:252] = w_color; end
            22 : begin tmp_color[275:264] = w_color; end
            23 : begin tmp_color[287:276] = w_color; end
            24 : begin tmp_color[299:288] = w_color; end
            25 : begin tmp_color[311:300] = w_color; end
            26 : begin tmp_color[323:312] = w_color; end
            27 : begin tmp_color[335:324] = w_color; end
            28 : begin tmp_color[347:336] = w_color; end
            29 : begin tmp_color[359:348] = w_color; end
            30 : begin tmp_color[371:360] = w_color; end
            31 : begin tmp_color[383:372] = w_color; end
            32 : begin tmp_color[395:384] = w_color; end
            33 : begin tmp_color[407:396] = w_color; end
            34 : begin tmp_color[419:408] = w_color; end
            35 : begin tmp_color[431:420] = w_color; end
            36 : begin tmp_color[443:432] = w_color; end
            37 : begin tmp_color[455:444] = w_color; end
            38 : begin tmp_color[467:456] = w_color; end
            39 : begin tmp_color[479:468] = w_color; end
            40 : begin tmp_color[491:480] = w_color; end
            41 : begin tmp_color[503:492] = w_color; end
            42 : begin tmp_color[515:504] = w_color; end
            43 : begin tmp_color[527:516] = w_color; end
            44 : begin tmp_color[539:528] = w_color; end
            45 : begin tmp_color[551:540] = w_color; end
            46 : begin tmp_color[563:552] = w_color; end
            47 : begin tmp_color[575:564] = w_color; end
            48 : begin tmp_color[587:576] = w_color; end
            49 : begin tmp_color[599:588] = w_color; end
            50 : begin tmp_color[611:600] = w_color; end
            51 : begin tmp_color[623:612] = w_color; end
            52 : begin tmp_color[635:624] = w_color; end
            53 : begin tmp_color[647:636] = w_color; end
            54 : begin tmp_color[659:648] = w_color; end
            55 : begin tmp_color[671:660] = w_color; end
            56 : begin tmp_color[683:672] = w_color; end
            57 : begin tmp_color[695:684] = w_color; end
            58 : begin tmp_color[707:696] = w_color; end
            59 : begin tmp_color[719:708] = w_color; end
            60 : begin tmp_color[731:720] = w_color; end
            61 : begin tmp_color[743:732] = w_color; end
            62 : begin tmp_color[755:744] = w_color; end
            63 : begin tmp_color[767:756] = w_color; end
            64 : begin tmp_color[779:768] = w_color; end
            65 : begin tmp_color[791:780] = w_color; end
            66 : begin tmp_color[803:792] = w_color; end
            67 : begin tmp_color[815:804] = w_color; end
            68 : begin tmp_color[827:816] = w_color; end
            69 : begin tmp_color[839:828] = w_color; end
            70 : begin tmp_color[851:840] = w_color; end
            71 : begin tmp_color[863:852] = w_color; end
            72 : begin tmp_color[875:864] = w_color; end
            73 : begin tmp_color[887:876] = w_color; end
            74 : begin tmp_color[899:888] = w_color; end
            75 : begin tmp_color[911:900] = w_color; end
            76 : begin tmp_color[923:912] = w_color; end
            77 : begin tmp_color[935:924] = w_color; end
            78 : begin tmp_color[947:936] = w_color; end
            79 : begin tmp_color[959:948] = w_color; end
            80 : begin tmp_color[971:960] = w_color; end
            81 : begin tmp_color[983:972] = w_color; end
            82 : begin tmp_color[995:984] = w_color; end
            83 : begin tmp_color[1007:996] = w_color; end
            84 : begin tmp_color[1019:1008] = w_color; end
            85 : begin tmp_color[1031:1020] = w_color; end
            86 : begin tmp_color[1043:1032] = w_color; end
            87 : begin tmp_color[1055:1044] = w_color; end
            88 : begin tmp_color[1067:1056] = w_color; end
            89 : begin tmp_color[1079:1068] = w_color; end
            90 : begin tmp_color[1091:1080] = w_color; end
            91 : begin tmp_color[1103:1092] = w_color; end
            92 : begin tmp_color[1115:1104] = w_color; end
            93 : begin tmp_color[1127:1116] = w_color; end
            94 : begin tmp_color[1139:1128] = w_color; end
            95 : begin tmp_color[1151:1140] = w_color; end
            96 : begin tmp_color[1163:1152] = w_color; end
            97 : begin tmp_color[1175:1164] = w_color; end
            98 : begin tmp_color[1187:1176] = w_color; end
            99 : begin tmp_color[1199:1188] = w_color; end
            100 : begin tmp_color[1211:1200] = w_color; end
            101 : begin tmp_color[1223:1212] = w_color; end
            102 : begin tmp_color[1235:1224] = w_color; end
            103 : begin tmp_color[1247:1236] = w_color; end
            104 : begin tmp_color[1259:1248] = w_color; end
            105 : begin tmp_color[1271:1260] = w_color; end
            106 : begin tmp_color[1283:1272] = w_color; end
            107 : begin tmp_color[1295:1284] = w_color; end
            108 : begin tmp_color[1307:1296] = w_color; end
            109 : begin tmp_color[1319:1308] = w_color; end
            110 : begin tmp_color[1331:1320] = w_color; end
            111 : begin tmp_color[1343:1332] = w_color; end
            112 : begin tmp_color[1355:1344] = w_color; end
            113 : begin tmp_color[1367:1356] = w_color; end
            114 : begin tmp_color[1379:1368] = w_color; end
            115 : begin tmp_color[1391:1380] = w_color; end
            116 : begin tmp_color[1403:1392] = w_color; end
            117 : begin tmp_color[1415:1404] = w_color; end
            118 : begin tmp_color[1427:1416] = w_color; end
            119 : begin tmp_color[1439:1428] = w_color; end
            120 : begin tmp_color[1451:1440] = w_color; end
            121 : begin tmp_color[1463:1452] = w_color; end
            122 : begin tmp_color[1475:1464] = w_color; end
            123 : begin tmp_color[1487:1476] = w_color; end
            124 : begin tmp_color[1499:1488] = w_color; end
            125 : begin tmp_color[1511:1500] = w_color; end
            126 : begin tmp_color[1523:1512] = w_color; end
            127 : begin tmp_color[1535:1524] = w_color; end
            128 : begin tmp_color[1547:1536] = w_color; end
            129 : begin tmp_color[1559:1548] = w_color; end
            130 : begin tmp_color[1571:1560] = w_color; end
            131 : begin tmp_color[1583:1572] = w_color; end
            132 : begin tmp_color[1595:1584] = w_color; end
            133 : begin tmp_color[1607:1596] = w_color; end
            134 : begin tmp_color[1619:1608] = w_color; end
            135 : begin tmp_color[1631:1620] = w_color; end
            136 : begin tmp_color[1643:1632] = w_color; end
            137 : begin tmp_color[1655:1644] = w_color; end
            138 : begin tmp_color[1667:1656] = w_color; end
            139 : begin tmp_color[1679:1668] = w_color; end
            140 : begin tmp_color[1691:1680] = w_color; end
            141 : begin tmp_color[1703:1692] = w_color; end
            142 : begin tmp_color[1715:1704] = w_color; end
            143 : begin tmp_color[1727:1716] = w_color; end
            144 : begin tmp_color[1739:1728] = w_color; end
            145 : begin tmp_color[1751:1740] = w_color; end
            146 : begin tmp_color[1763:1752] = w_color; end
            147 : begin tmp_color[1775:1764] = w_color; end
            148 : begin tmp_color[1787:1776] = w_color; end
            149 : begin tmp_color[1799:1788] = w_color; end
            150 : begin tmp_color[1811:1800] = w_color; end
            151 : begin tmp_color[1823:1812] = w_color; end
            152 : begin tmp_color[1835:1824] = w_color; end
            153 : begin tmp_color[1847:1836] = w_color; end
            154 : begin tmp_color[1859:1848] = w_color; end
            155 : begin tmp_color[1871:1860] = w_color; end
            156 : begin tmp_color[1883:1872] = w_color; end
            157 : begin tmp_color[1895:1884] = w_color; end
            158 : begin tmp_color[1907:1896] = w_color; end
            159 : begin tmp_color[1919:1908] = w_color; end
            160 : begin tmp_color[1931:1920] = w_color; end
            161 : begin tmp_color[1943:1932] = w_color; end
            162 : begin tmp_color[1955:1944] = w_color; end
            163 : begin tmp_color[1967:1956] = w_color; end
            164 : begin tmp_color[1979:1968] = w_color; end
            165 : begin tmp_color[1991:1980] = w_color; end
            166 : begin tmp_color[2003:1992] = w_color; end
            167 : begin tmp_color[2015:2004] = w_color; end
            168 : begin tmp_color[2027:2016] = w_color; end
            169 : begin tmp_color[2039:2028] = w_color; end
            170 : begin tmp_color[2051:2040] = w_color; end
            171 : begin tmp_color[2063:2052] = w_color; end
            172 : begin tmp_color[2075:2064] = w_color; end
            173 : begin tmp_color[2087:2076] = w_color; end
            174 : begin tmp_color[2099:2088] = w_color; end
            175 : begin tmp_color[2111:2100] = w_color; end
            176 : begin tmp_color[2123:2112] = w_color; end
            177 : begin tmp_color[2135:2124] = w_color; end
            178 : begin tmp_color[2147:2136] = w_color; end
            179 : begin tmp_color[2159:2148] = w_color; end
            180 : begin tmp_color[2171:2160] = w_color; end
            181 : begin tmp_color[2183:2172] = w_color; end
            182 : begin tmp_color[2195:2184] = w_color; end
            183 : begin tmp_color[2207:2196] = w_color; end
            184 : begin tmp_color[2219:2208] = w_color; end
            185 : begin tmp_color[2231:2220] = w_color; end
            186 : begin tmp_color[2243:2232] = w_color; end
            187 : begin tmp_color[2255:2244] = w_color; end
            188 : begin tmp_color[2267:2256] = w_color; end
            189 : begin tmp_color[2279:2268] = w_color; end
            190 : begin tmp_color[2291:2280] = w_color; end
            191 : begin tmp_color[2303:2292] = w_color; end
            192 : begin tmp_color[2315:2304] = w_color; end
            193 : begin tmp_color[2327:2316] = w_color; end
            194 : begin tmp_color[2339:2328] = w_color; end
            195 : begin tmp_color[2351:2340] = w_color; end
            196 : begin tmp_color[2363:2352] = w_color; end
            197 : begin tmp_color[2375:2364] = w_color; end
            198 : begin tmp_color[2387:2376] = w_color; end
            199 : begin tmp_color[2399:2388] = w_color; end
            200 : begin tmp_color[2411:2400] = w_color; end
            201 : begin tmp_color[2423:2412] = w_color; end
            202 : begin tmp_color[2435:2424] = w_color; end
            203 : begin tmp_color[2447:2436] = w_color; end
            204 : begin tmp_color[2459:2448] = w_color; end
            205 : begin tmp_color[2471:2460] = w_color; end
            206 : begin tmp_color[2483:2472] = w_color; end
            207 : begin tmp_color[2495:2484] = w_color; end
            208 : begin tmp_color[2507:2496] = w_color; end
            209 : begin tmp_color[2519:2508] = w_color; end
            210 : begin tmp_color[2531:2520] = w_color; end
            211 : begin tmp_color[2543:2532] = w_color; end
            212 : begin tmp_color[2555:2544] = w_color; end
            213 : begin tmp_color[2567:2556] = w_color; end
            214 : begin tmp_color[2579:2568] = w_color; end
            215 : begin tmp_color[2591:2580] = w_color; end
            216 : begin tmp_color[2603:2592] = w_color; end
            217 : begin tmp_color[2615:2604] = w_color; end
            218 : begin tmp_color[2627:2616] = w_color; end
            219 : begin tmp_color[2639:2628] = w_color; end
            220 : begin tmp_color[2651:2640] = w_color; end
            221 : begin tmp_color[2663:2652] = w_color; end
            222 : begin tmp_color[2675:2664] = w_color; end
            223 : begin tmp_color[2687:2676] = w_color; end
            224 : begin tmp_color[2699:2688] = w_color; end
            225 : begin tmp_color[2711:2700] = w_color; end
            226 : begin tmp_color[2723:2712] = w_color; end
            227 : begin tmp_color[2735:2724] = w_color; end
            228 : begin tmp_color[2747:2736] = w_color; end
            229 : begin tmp_color[2759:2748] = w_color; end
            230 : begin tmp_color[2771:2760] = w_color; end
            231 : begin tmp_color[2783:2772] = w_color; end
            232 : begin tmp_color[2795:2784] = w_color; end
            233 : begin tmp_color[2807:2796] = w_color; end
            234 : begin tmp_color[2819:2808] = w_color; end
            235 : begin tmp_color[2831:2820] = w_color; end
            236 : begin tmp_color[2843:2832] = w_color; end
            237 : begin tmp_color[2855:2844] = w_color; end
            238 : begin tmp_color[2867:2856] = w_color; end
            239 : begin tmp_color[2879:2868] = w_color; end
            default:begin end
        endcase
    end
    else begin
            tmp_color[11:0] = (block_exist[0])?color[11:0]:12'h111;
            tmp_color[23:12] = (block_exist[1])?color[23:12]:12'h222;
            tmp_color[35:24] = (block_exist[2])?color[35:24]:12'h111;
            tmp_color[47:36] = (block_exist[3])?color[47:36]:12'h222;
            tmp_color[59:48] = (block_exist[4])?color[59:48]:12'h111;
            tmp_color[71:60] = (block_exist[5])?color[71:60]:12'h222;
            tmp_color[83:72] = (block_exist[6])?color[83:72]:12'h111;
            tmp_color[95:84] = (block_exist[7])?color[95:84]:12'h222;
            tmp_color[107:96] = (block_exist[8])?color[107:96]:12'h111;
            tmp_color[119:108] = (block_exist[9])?color[119:108]:12'h222;
            tmp_color[131:120] = (block_exist[10])?color[131:120]:12'h222;
            tmp_color[143:132] = (block_exist[11])?color[143:132]:12'h111;
            tmp_color[155:144] = (block_exist[12])?color[155:144]:12'h222;
            tmp_color[167:156] = (block_exist[13])?color[167:156]:12'h111;
            tmp_color[179:168] = (block_exist[14])?color[179:168]:12'h222;
            tmp_color[191:180] = (block_exist[15])?color[191:180]:12'h111;
            tmp_color[203:192] = (block_exist[16])?color[203:192]:12'h222;
            tmp_color[215:204] = (block_exist[17])?color[215:204]:12'h111;
            tmp_color[227:216] = (block_exist[18])?color[227:216]:12'h222;
            tmp_color[239:228] = (block_exist[19])?color[239:228]:12'h111;
            tmp_color[251:240] = (block_exist[20])?color[251:240]:12'h111;
            tmp_color[263:252] = (block_exist[21])?color[263:252]:12'h222;
            tmp_color[275:264] = (block_exist[22])?color[275:264]:12'h111;
            tmp_color[287:276] = (block_exist[23])?color[287:276]:12'h222;
            tmp_color[299:288] = (block_exist[24])?color[299:288]:12'h111;
            tmp_color[311:300] = (block_exist[25])?color[311:300]:12'h222;
            tmp_color[323:312] = (block_exist[26])?color[323:312]:12'h111;
            tmp_color[335:324] = (block_exist[27])?color[335:324]:12'h222;
            tmp_color[347:336] = (block_exist[28])?color[347:336]:12'h111;
            tmp_color[359:348] = (block_exist[29])?color[359:348]:12'h222;
            tmp_color[371:360] = (block_exist[30])?color[371:360]:12'h222;
            tmp_color[383:372] = (block_exist[31])?color[383:372]:12'h111;
            tmp_color[395:384] = (block_exist[32])?color[395:384]:12'h222;
            tmp_color[407:396] = (block_exist[33])?color[407:396]:12'h111;
            tmp_color[419:408] = (block_exist[34])?color[419:408]:12'h222;
            tmp_color[431:420] = (block_exist[35])?color[431:420]:12'h111;
            tmp_color[443:432] = (block_exist[36])?color[443:432]:12'h222;
            tmp_color[455:444] = (block_exist[37])?color[455:444]:12'h111;
            tmp_color[467:456] = (block_exist[38])?color[467:456]:12'h222;
            tmp_color[479:468] = (block_exist[39])?color[479:468]:12'h111;
            tmp_color[491:480] = (block_exist[40])?color[491:480]:12'h111;
            tmp_color[503:492] = (block_exist[41])?color[503:492]:12'h222;
            tmp_color[515:504] = (block_exist[42])?color[515:504]:12'h111;
            tmp_color[527:516] = (block_exist[43])?color[527:516]:12'h222;
            tmp_color[539:528] = (block_exist[44])?color[539:528]:12'h111;
            tmp_color[551:540] = (block_exist[45])?color[551:540]:12'h222;
            tmp_color[563:552] = (block_exist[46])?color[563:552]:12'h111;
            tmp_color[575:564] = (block_exist[47])?color[575:564]:12'h222;
            tmp_color[587:576] = (block_exist[48])?color[587:576]:12'h111;
            tmp_color[599:588] = (block_exist[49])?color[599:588]:12'h222;
            tmp_color[611:600] = (block_exist[50])?color[611:600]:12'h222;
            tmp_color[623:612] = (block_exist[51])?color[623:612]:12'h111;
            tmp_color[635:624] = (block_exist[52])?color[635:624]:12'h222;
            tmp_color[647:636] = (block_exist[53])?color[647:636]:12'h111;
            tmp_color[659:648] = (block_exist[54])?color[659:648]:12'h222;
            tmp_color[671:660] = (block_exist[55])?color[671:660]:12'h111;
            tmp_color[683:672] = (block_exist[56])?color[683:672]:12'h222;
            tmp_color[695:684] = (block_exist[57])?color[695:684]:12'h111;
            tmp_color[707:696] = (block_exist[58])?color[707:696]:12'h222;
            tmp_color[719:708] = (block_exist[59])?color[719:708]:12'h111;
            tmp_color[731:720] = (block_exist[60])?color[731:720]:12'h111;
            tmp_color[743:732] = (block_exist[61])?color[743:732]:12'h222;
            tmp_color[755:744] = (block_exist[62])?color[755:744]:12'h111;
            tmp_color[767:756] = (block_exist[63])?color[767:756]:12'h222;
            tmp_color[779:768] = (block_exist[64])?color[779:768]:12'h111;
            tmp_color[791:780] = (block_exist[65])?color[791:780]:12'h222;
            tmp_color[803:792] = (block_exist[66])?color[803:792]:12'h111;
            tmp_color[815:804] = (block_exist[67])?color[815:804]:12'h222;
            tmp_color[827:816] = (block_exist[68])?color[827:816]:12'h111;
            tmp_color[839:828] = (block_exist[69])?color[839:828]:12'h222;
            tmp_color[851:840] = (block_exist[70])?color[851:840]:12'h222;
            tmp_color[863:852] = (block_exist[71])?color[863:852]:12'h111;
            tmp_color[875:864] = (block_exist[72])?color[875:864]:12'h222;
            tmp_color[887:876] = (block_exist[73])?color[887:876]:12'h111;
            tmp_color[899:888] = (block_exist[74])?color[899:888]:12'h222;
            tmp_color[911:900] = (block_exist[75])?color[911:900]:12'h111;
            tmp_color[923:912] = (block_exist[76])?color[923:912]:12'h222;
            tmp_color[935:924] = (block_exist[77])?color[935:924]:12'h111;
            tmp_color[947:936] = (block_exist[78])?color[947:936]:12'h222;
            tmp_color[959:948] = (block_exist[79])?color[959:948]:12'h111;
            tmp_color[971:960] = (block_exist[80])?color[971:960]:12'h111;
            tmp_color[983:972] = (block_exist[81])?color[983:972]:12'h222;
            tmp_color[995:984] = (block_exist[82])?color[995:984]:12'h111;
            tmp_color[1007:996] = (block_exist[83])?color[1007:996]:12'h222; 
            tmp_color[1019:1008] = (block_exist[84])?color[1019:1008]:12'h111;
            tmp_color[1031:1020] = (block_exist[85])?color[1031:1020]:12'h222;
            tmp_color[1043:1032] = (block_exist[86])?color[1043:1032]:12'h111;
            tmp_color[1055:1044] = (block_exist[87])?color[1055:1044]:12'h222;
            tmp_color[1067:1056] = (block_exist[88])?color[1067:1056]:12'h111;
            tmp_color[1079:1068] = (block_exist[89])?color[1079:1068]:12'h222;
            tmp_color[1091:1080] = (block_exist[90])?color[1091:1080]:12'h222;
            tmp_color[1103:1092] = (block_exist[91])?color[1103:1092]:12'h111;
            tmp_color[1115:1104] = (block_exist[92])?color[1115:1104]:12'h222;
            tmp_color[1127:1116] = (block_exist[93])?color[1127:1116]:12'h111;
            tmp_color[1139:1128] = (block_exist[94])?color[1139:1128]:12'h222;
            tmp_color[1151:1140] = (block_exist[95])?color[1151:1140]:12'h111;
            tmp_color[1163:1152] = (block_exist[96])?color[1163:1152]:12'h222;
            tmp_color[1175:1164] = (block_exist[97])?color[1175:1164]:12'h111;
            tmp_color[1187:1176] = (block_exist[98])?color[1187:1176]:12'h222;
            tmp_color[1199:1188] = (block_exist[99])?color[1199:1188]:12'h111;
            tmp_color[1211:1200] = (block_exist[100])?color[1211:1200]:12'h111;
            tmp_color[1223:1212] = (block_exist[101])?color[1223:1212]:12'h222;
            tmp_color[1235:1224] = (block_exist[102])?color[1235:1224]:12'h111;
            tmp_color[1247:1236] = (block_exist[103])?color[1247:1236]:12'h222;
            tmp_color[1259:1248] = (block_exist[104])?color[1259:1248]:12'h111;
            tmp_color[1271:1260] = (block_exist[105])?color[1271:1260]:12'h222;
            tmp_color[1283:1272] = (block_exist[106])?color[1283:1272]:12'h111;
            tmp_color[1295:1284] = (block_exist[107])?color[1295:1284]:12'h222;
            tmp_color[1307:1296] = (block_exist[108])?color[1307:1296]:12'h111;
            tmp_color[1319:1308] = (block_exist[109])?color[1319:1308]:12'h222;
            tmp_color[1331:1320] = (block_exist[110])?color[1331:1320]:12'h222;
            tmp_color[1343:1332] = (block_exist[111])?color[1343:1332]:12'h111;
            tmp_color[1355:1344] = (block_exist[112])?color[1355:1344]:12'h222;
            tmp_color[1367:1356] = (block_exist[113])?color[1367:1356]:12'h111;
            tmp_color[1379:1368] = (block_exist[114])?color[1379:1368]:12'h222;
            tmp_color[1391:1380] = (block_exist[115])?color[1391:1380]:12'h111;
            tmp_color[1403:1392] = (block_exist[116])?color[1403:1392]:12'h222;
            tmp_color[1415:1404] = (block_exist[117])?color[1415:1404]:12'h111;
            tmp_color[1427:1416] = (block_exist[118])?color[1427:1416]:12'h222;
            tmp_color[1439:1428] = (block_exist[119])?color[1439:1428]:12'h111;
            tmp_color[1451:1440] = (block_exist[120])?color[1451:1440]:12'h111;
            tmp_color[1463:1452] = (block_exist[121])?color[1463:1452]:12'h222;
            tmp_color[1475:1464] = (block_exist[122])?color[1475:1464]:12'h111;
            tmp_color[1487:1476] = (block_exist[123])?color[1487:1476]:12'h222;
            tmp_color[1499:1488] = (block_exist[124])?color[1499:1488]:12'h111;
            tmp_color[1511:1500] = (block_exist[125])?color[1511:1500]:12'h222;
            tmp_color[1523:1512] = (block_exist[126])?color[1523:1512]:12'h111;
            tmp_color[1535:1524] = (block_exist[127])?color[1535:1524]:12'h222;
            tmp_color[1547:1536] = (block_exist[128])?color[1547:1536]:12'h111;
            tmp_color[1559:1548] = (block_exist[129])?color[1559:1548]:12'h222;
            tmp_color[1571:1560] = (block_exist[130])?color[1571:1560]:12'h222;
            tmp_color[1583:1572] = (block_exist[131])?color[1583:1572]:12'h111;
            tmp_color[1595:1584] = (block_exist[132])?color[1595:1584]:12'h222;
            tmp_color[1607:1596] = (block_exist[133])?color[1607:1596]:12'h111;
            tmp_color[1619:1608] = (block_exist[134])?color[1619:1608]:12'h222;
            tmp_color[1631:1620] = (block_exist[135])?color[1631:1620]:12'h111;
            tmp_color[1643:1632] = (block_exist[136])?color[1643:1632]:12'h222;
            tmp_color[1655:1644] = (block_exist[137])?color[1655:1644]:12'h111;
            tmp_color[1667:1656] = (block_exist[138])?color[1667:1656]:12'h222;
            tmp_color[1679:1668] = (block_exist[139])?color[1679:1668]:12'h111;
            tmp_color[1691:1680] = (block_exist[140])?color[1691:1680]:12'h111;
            tmp_color[1703:1692] = (block_exist[141])?color[1703:1692]:12'h222;
            tmp_color[1715:1704] = (block_exist[142])?color[1715:1704]:12'h111;
            tmp_color[1727:1716] = (block_exist[143])?color[1727:1716]:12'h222;
            tmp_color[1739:1728] = (block_exist[144])?color[1739:1728]:12'h111;
            tmp_color[1751:1740] = (block_exist[145])?color[1751:1740]:12'h222;
            tmp_color[1763:1752] = (block_exist[146])?color[1763:1752]:12'h111;
            tmp_color[1775:1764] = (block_exist[147])?color[1775:1764]:12'h222;
            tmp_color[1787:1776] = (block_exist[148])?color[1787:1776]:12'h111;
            tmp_color[1799:1788] = (block_exist[149])?color[1799:1788]:12'h222;
            tmp_color[1811:1800] = (block_exist[150])?color[1811:1800]:12'h222;
            tmp_color[1823:1812] = (block_exist[151])?color[1823:1812]:12'h111;
            tmp_color[1835:1824] = (block_exist[152])?color[1835:1824]:12'h222;
            tmp_color[1847:1836] = (block_exist[153])?color[1847:1836]:12'h111;
            tmp_color[1859:1848] = (block_exist[154])?color[1859:1848]:12'h222;
            tmp_color[1871:1860] = (block_exist[155])?color[1871:1860]:12'h111;
            tmp_color[1883:1872] = (block_exist[156])?color[1883:1872]:12'h222;
            tmp_color[1895:1884] = (block_exist[157])?color[1895:1884]:12'h111;
            tmp_color[1907:1896] = (block_exist[158])?color[1907:1896]:12'h222;
            tmp_color[1919:1908] = (block_exist[159])?color[1919:1908]:12'h111;
            tmp_color[1931:1920] = (block_exist[160])?color[1931:1920]:12'h111;
            tmp_color[1943:1932] = (block_exist[161])?color[1943:1932]:12'h222;
            tmp_color[1955:1944] = (block_exist[162])?color[1955:1944]:12'h111;
            tmp_color[1967:1956] = (block_exist[163])?color[1967:1956]:12'h222;
            tmp_color[1979:1968] = (block_exist[164])?color[1979:1968]:12'h111;
            tmp_color[1991:1980] = (block_exist[165])?color[1991:1980]:12'h222;
            tmp_color[2003:1992] = (block_exist[166])?color[2003:1992]:12'h111;
            tmp_color[2015:2004] = (block_exist[167])?color[2015:2004]:12'h222;
            tmp_color[2027:2016] = (block_exist[168])?color[2027:2016]:12'h111;
            tmp_color[2039:2028] = (block_exist[169])?color[2039:2028]:12'h222;
            tmp_color[2051:2040] = (block_exist[170])?color[2051:2040]:12'h222;
            tmp_color[2063:2052] = (block_exist[171])?color[2063:2052]:12'h111;
            tmp_color[2075:2064] = (block_exist[172])?color[2075:2064]:12'h222;
            tmp_color[2087:2076] = (block_exist[173])?color[2087:2076]:12'h111;
            tmp_color[2099:2088] = (block_exist[174])?color[2099:2088]:12'h222;
            tmp_color[2111:2100] = (block_exist[175])?color[2111:2100]:12'h111;
            tmp_color[2123:2112] = (block_exist[176])?color[2123:2112]:12'h222;
            tmp_color[2135:2124] = (block_exist[177])?color[2135:2124]:12'h111;
            tmp_color[2147:2136] = (block_exist[178])?color[2147:2136]:12'h222;
            tmp_color[2159:2148] = (block_exist[179])?color[2159:2148]:12'h111;
            tmp_color[2171:2160] = (block_exist[180])?color[2171:2160]:12'h111;
            tmp_color[2183:2172] = (block_exist[181])?color[2183:2172]:12'h222;
            tmp_color[2195:2184] = (block_exist[182])?color[2195:2184]:12'h111;
            tmp_color[2207:2196] = (block_exist[183])?color[2207:2196]:12'h222;
            tmp_color[2219:2208] = (block_exist[184])?color[2219:2208]:12'h111;
            tmp_color[2231:2220] = (block_exist[185])?color[2231:2220]:12'h222;
            tmp_color[2243:2232] = (block_exist[186])?color[2243:2232]:12'h111;
            tmp_color[2255:2244] = (block_exist[187])?color[2255:2244]:12'h222;
            tmp_color[2267:2256] = (block_exist[188])?color[2267:2256]:12'h111;
            tmp_color[2279:2268] = (block_exist[189])?color[2279:2268]:12'h222;
            tmp_color[2291:2280] = (block_exist[190])?color[2291:2280]:12'h222;
            tmp_color[2303:2292] = (block_exist[191])?color[2303:2292]:12'h111;
            tmp_color[2315:2304] = (block_exist[192])?color[2315:2304]:12'h222;
            tmp_color[2327:2316] = (block_exist[193])?color[2327:2316]:12'h111;
            tmp_color[2339:2328] = (block_exist[194])?color[2339:2328]:12'h222;
            tmp_color[2351:2340] = (block_exist[195])?color[2351:2340]:12'h111;
            tmp_color[2363:2352] = (block_exist[196])?color[2363:2352]:12'h222;
            tmp_color[2375:2364] = (block_exist[197])?color[2375:2364]:12'h111;
            tmp_color[2387:2376] = (block_exist[198])?color[2387:2376]:12'h222;
            tmp_color[2399:2388] = (block_exist[199])?color[2399:2388]:12'h111;
            tmp_color[2411:2400] = (block_exist[200])?color[2411:2400]:12'h111;
            tmp_color[2423:2412] = (block_exist[201])?color[2423:2412]:12'h111;
            tmp_color[2435:2424] = (block_exist[202])?color[2435:2424]:12'h111;
            tmp_color[2447:2436] = (block_exist[203])?color[2447:2436]:12'h111;
            tmp_color[2459:2448] = (block_exist[204])?color[2459:2448]:12'h111;
            tmp_color[2471:2460] = (block_exist[205])?color[2471:2460]:12'h111;
            tmp_color[2483:2472] = (block_exist[206])?color[2483:2472]:12'h111;
            tmp_color[2495:2484] = (block_exist[207])?color[2495:2484]:12'h111;
            tmp_color[2507:2496] = (block_exist[208])?color[2507:2496]:12'h111;
            tmp_color[2519:2508] = (block_exist[209])?color[2519:2508]:12'h111;
            tmp_color[2531:2520] = (block_exist[210])?color[2531:2520]:12'h111;
            tmp_color[2543:2532] = (block_exist[211])?color[2543:2532]:12'h111;
            tmp_color[2555:2544] = (block_exist[212])?color[2555:2544]:12'h111;
            tmp_color[2567:2556] = (block_exist[213])?color[2567:2556]:12'h111;
            tmp_color[2579:2568] = (block_exist[214])?color[2579:2568]:12'h111;
            tmp_color[2591:2580] = (block_exist[215])?color[2591:2580]:12'h111;
            tmp_color[2603:2592] = (block_exist[216])?color[2603:2592]:12'h111;
            tmp_color[2615:2604] = (block_exist[217])?color[2615:2604]:12'h111;
            tmp_color[2627:2616] = (block_exist[218])?color[2627:2616]:12'h111;
            tmp_color[2639:2628] = (block_exist[219])?color[2639:2628]:12'h111;
            tmp_color[2651:2640] = (block_exist[220])?color[2651:2640]:12'h111;
            tmp_color[2663:2652] = (block_exist[221])?color[2663:2652]:12'h111;
            tmp_color[2675:2664] = (block_exist[222])?color[2675:2664]:12'h111;
            tmp_color[2687:2676] = (block_exist[223])?color[2687:2676]:12'h111;
            tmp_color[2699:2688] = (block_exist[224])?color[2699:2688]:12'h111;
            tmp_color[2711:2700] = (block_exist[225])?color[2711:2700]:12'h111;
            tmp_color[2723:2712] = (block_exist[226])?color[2723:2712]:12'h111;
            tmp_color[2735:2724] = (block_exist[227])?color[2735:2724]:12'h111;
            tmp_color[2747:2736] = (block_exist[228])?color[2747:2736]:12'h111;
            tmp_color[2759:2748] = (block_exist[229])?color[2759:2748]:12'h111;
            tmp_color[2771:2760] = (block_exist[230])?color[2771:2760]:12'h111;
            tmp_color[2783:2772] = (block_exist[231])?color[2783:2772]:12'h111;
            tmp_color[2795:2784] = (block_exist[232])?color[2795:2784]:12'h111;
            tmp_color[2807:2796] = (block_exist[233])?color[2807:2796]:12'h111;
            tmp_color[2819:2808] = (block_exist[234])?color[2819:2808]:12'h111;
            tmp_color[2831:2820] = (block_exist[235])?color[2831:2820]:12'h111;
            tmp_color[2843:2832] = (block_exist[236])?color[2843:2832]:12'h111;
            tmp_color[2855:2844] = (block_exist[237])?color[2855:2844]:12'h111;
            tmp_color[2867:2856] = (block_exist[238])?color[2867:2856]:12'h111;
            tmp_color[2879:2868] = (block_exist[239])?color[2879:2868]:12'h111;
    end
end
always@(posedge clk or posedge rst)begin
    if(rst)begin
        read_addr_color <= 12'h111;
        color[11:0]<=12'h111;
        color[23:12]<=12'h222;
        color[35:24]<=12'h111;
        color[47:36]<=12'h222;
        color[59:48]<=12'h111;
        color[71:60]<=12'h222;
        color[83:72]<=12'h111;
        color[95:84]<=12'h222;
        color[107:96]<=12'h111;
        color[119:108]<=12'h222;
        color[131:120]<=12'h222;
        color[143:132]<=12'h111;
        color[155:144]<=12'h222;
        color[167:156]<=12'h111;
        color[179:168]<=12'h222;
        color[191:180]<=12'h111;
        color[203:192]<=12'h222;
        color[215:204]<=12'h111;
        color[227:216]<=12'h222;
        color[239:228]<=12'h111;
        color[251:240]<=12'h111;
        color[263:252]<=12'h222;
        color[275:264]<=12'h111;
        color[287:276]<=12'h222;
        color[299:288]<=12'h111;
        color[311:300]<=12'h222;
        color[323:312]<=12'h111;
        color[335:324]<=12'h222;
        color[347:336]<=12'h111;
        color[359:348]<=12'h222;
        color[371:360]<=12'h222;
        color[383:372]<=12'h111;
        color[395:384]<=12'h222;
        color[407:396]<=12'h111;
        color[419:408]<=12'h222;
        color[431:420]<=12'h111;
        color[443:432]<=12'h222;
        color[455:444]<=12'h111;
        color[467:456]<=12'h222;
        color[479:468]<=12'h111;
        color[491:480]<=12'h111;
        color[503:492]<=12'h222;
        color[515:504]<=12'h111;
        color[527:516]<=12'h222;
        color[539:528]<=12'h111;
        color[551:540]<=12'h222;
        color[563:552]<=12'h111;
        color[575:564]<=12'h222;
        color[587:576]<=12'h111;
        color[599:588]<=12'h222;
        color[611:600]<=12'h222;
        color[623:612]<=12'h111;
        color[635:624]<=12'h222;
        color[647:636]<=12'h111;
        color[659:648]<=12'h222;
        color[671:660]<=12'h111;
        color[683:672]<=12'h222;
        color[695:684]<=12'h111;
        color[707:696]<=12'h222;
        color[719:708]<=12'h111;
        color[731:720]<=12'h111;
        color[743:732]<=12'h222;
        color[755:744]<=12'h111;
        color[767:756]<=12'h222;
        color[779:768]<=12'h111;
        color[791:780]<=12'h222;
        color[803:792]<=12'h111;
        color[815:804]<=12'h222;
        color[827:816]<=12'h111;
        color[839:828]<=12'h222;
        color[851:840]<=12'h222;
        color[863:852]<=12'h111;
        color[875:864]<=12'h222;
        color[887:876]<=12'h111;
        color[899:888]<=12'h222;
        color[911:900]<=12'h111;
        color[923:912]<=12'h222;
        color[935:924]<=12'h111;
        color[947:936]<=12'h222;
        color[959:948]<=12'h111;
        color[971:960]<=12'h111;
        color[983:972]<=12'h222;
        color[995:984]<=12'h111;
        color[1007:996]<=12'h222;
        color[1019:1008]<=12'h111;
        color[1031:1020]<=12'h222;
        color[1043:1032]<=12'h111;
        color[1055:1044]<=12'h222;
        color[1067:1056]<=12'h111;
        color[1079:1068]<=12'h222;
        color[1091:1080]<=12'h222;
        color[1103:1092]<=12'h111;
        color[1115:1104]<=12'h222;
        color[1127:1116]<=12'h111;
        color[1139:1128]<=12'h222;
        color[1151:1140]<=12'h111;
        color[1163:1152]<=12'h222;
        color[1175:1164]<=12'h111;
        color[1187:1176]<=12'h222;
        color[1199:1188]<=12'h111;
        color[1211:1200]<=12'h111;
        color[1223:1212]<=12'h222;
        color[1235:1224]<=12'h111;
        color[1247:1236]<=12'h222;
        color[1259:1248]<=12'h111;
        color[1271:1260]<=12'h222;
        color[1283:1272]<=12'h111;
        color[1295:1284]<=12'h222;
        color[1307:1296]<=12'h111;
        color[1319:1308]<=12'h222;
        color[1331:1320]<=12'h222;
        color[1343:1332]<=12'h111;
        color[1355:1344]<=12'h222;
        color[1367:1356]<=12'h111;
        color[1379:1368]<=12'h222;
        color[1391:1380]<=12'h111;
        color[1403:1392]<=12'h222;
        color[1415:1404]<=12'h111;
        color[1427:1416]<=12'h222;
        color[1439:1428]<=12'h111;
        color[1451:1440]<=12'h111;
        color[1463:1452]<=12'h222;
        color[1475:1464]<=12'h111;
        color[1487:1476]<=12'h222;
        color[1499:1488]<=12'h111;
        color[1511:1500]<=12'h222;
        color[1523:1512]<=12'h111;
        color[1535:1524]<=12'h222;
        color[1547:1536]<=12'h111;
        color[1559:1548]<=12'h222;
        color[1571:1560]<=12'h222;
        color[1583:1572]<=12'h111;
        color[1595:1584]<=12'h222;
        color[1607:1596]<=12'h111;
        color[1619:1608]<=12'h222;
        color[1631:1620]<=12'h111;
        color[1643:1632]<=12'h222;
        color[1655:1644]<=12'h111;
        color[1667:1656]<=12'h222;
        color[1679:1668]<=12'h111;
        color[1691:1680]<=12'h111;
        color[1703:1692]<=12'h222;
        color[1715:1704]<=12'h111;
        color[1727:1716]<=12'h222;
        color[1739:1728]<=12'h111;
        color[1751:1740]<=12'h222;
        color[1763:1752]<=12'h111;
        color[1775:1764]<=12'h222;
        color[1787:1776]<=12'h111;
        color[1799:1788]<=12'h222;
        color[1811:1800]<=12'h222;
        color[1823:1812]<=12'h111;
        color[1835:1824]<=12'h222;
        color[1847:1836]<=12'h111;
        color[1859:1848]<=12'h222;
        color[1871:1860]<=12'h111;
        color[1883:1872]<=12'h222;
        color[1895:1884]<=12'h111;
        color[1907:1896]<=12'h222;
        color[1919:1908]<=12'h111;
        color[1931:1920]<=12'h111;
        color[1943:1932]<=12'h222;
        color[1955:1944]<=12'h111;
        color[1967:1956]<=12'h222;
        color[1979:1968]<=12'h111;
        color[1991:1980]<=12'h222;
        color[2003:1992]<=12'h111;
        color[2015:2004]<=12'h222;
        color[2027:2016]<=12'h111;
        color[2039:2028]<=12'h222;
        color[2051:2040]<=12'h222;
        color[2063:2052]<=12'h111;
        color[2075:2064]<=12'h222;
        color[2087:2076]<=12'h111;
        color[2099:2088]<=12'h222;
        color[2111:2100]<=12'h111;
        color[2123:2112]<=12'h222;
        color[2135:2124]<=12'h111;
        color[2147:2136]<=12'h222;
        color[2159:2148]<=12'h111;
        color[2171:2160]<=12'h111;
        color[2183:2172]<=12'h222;
        color[2195:2184]<=12'h111;
        color[2207:2196]<=12'h222;
        color[2219:2208]<=12'h111;
        color[2231:2220]<=12'h222;
        color[2243:2232]<=12'h111;
        color[2255:2244]<=12'h222;
        color[2267:2256]<=12'h111;
        color[2279:2268]<=12'h222;
        color[2291:2280]<=12'h222;
        color[2303:2292]<=12'h111;
        color[2315:2304]<=12'h222;
        color[2327:2316]<=12'h111;
        color[2339:2328]<=12'h222;
        color[2351:2340]<=12'h111;
        color[2363:2352]<=12'h222;
        color[2375:2364]<=12'h111;
        color[2387:2376]<=12'h222;
        color[2399:2388]<=12'h111;
        color[2411:2400]<=12'h111;
        color[2423:2412]<=12'h111;
        color[2435:2424]<=12'h111;
        color[2447:2436]<=12'h111;
        color[2459:2448]<=12'h111;
        color[2471:2460]<=12'h111;
        color[2483:2472]<=12'h111;
        color[2495:2484]<=12'h111;
        color[2507:2496]<=12'h111;
        color[2519:2508]<=12'h111;
        color[2531:2520]<=12'h111;
        color[2543:2532]<=12'h111;
        color[2555:2544]<=12'h111;
        color[2567:2556]<=12'h111;
        color[2579:2568]<=12'h111;
        color[2591:2580]<=12'h111;
        color[2603:2592]<=12'h111;
        color[2615:2604]<=12'h111;
        color[2627:2616]<=12'h111;
        color[2639:2628]<=12'h111;
        color[2651:2640]<=12'h111;
        color[2663:2652]<=12'h111;
        color[2675:2664]<=12'h111;
        color[2687:2676]<=12'h111;
        color[2699:2688]<=12'h111;
        color[2711:2700]<=12'h111;
        color[2723:2712]<=12'h111;
        color[2735:2724]<=12'h111;
        color[2747:2736]<=12'h111;
        color[2759:2748]<=12'h111;
        color[2771:2760]<=12'h111;
        color[2783:2772]<=12'h111;
        color[2795:2784]<=12'h111;
        color[2807:2796]<=12'h111;
        color[2819:2808]<=12'h111;
        color[2831:2820]<=12'h111;
        color[2843:2832]<=12'h111;
        color[2855:2844]<=12'h111;
        color[2867:2856]<=12'h111;
        color[2879:2868]<=12'h111;  
foresee[11:0]<=12'h222;
foresee[23:12]<=12'h111;
foresee[35:24]<=12'h222;
foresee[47:36]<=12'h111;
foresee[59:48]<=12'h222;
foresee[71:60]<=12'h111;
foresee[83:72]<=12'h222;
foresee[95:84]<=12'h111;
foresee[107:96]<=12'h222;
foresee[119:108]<=12'h111;
foresee[131:120]<=12'h222;
foresee[143:132]<=12'h111;
foresee[155:144]<=12'h222;
foresee[167:156]<=12'h111;
foresee[179:168]<=12'h222;
foresee[191:180]<=12'h111;
foresee[203:192]<=12'h222;
foresee[215:204]<=12'h111;
foresee[227:216]<=12'h222;
foresee[239:228]<=12'h111;
foresee[251:240]<=12'h222;
foresee[263:252]<=12'h111;
foresee[275:264]<=12'h222;
foresee[287:276]<=12'h111;
foresee[299:288]<=12'h222;
foresee[311:300]<=12'h111;
foresee[323:312]<=12'h222;
foresee[335:324]<=12'h111;
foresee[347:336]<=12'h222;
foresee[359:348]<=12'h111;
foresee[371:360]<=12'h222;
foresee[383:372]<=12'h111;
foresee[395:384]<=12'h222;
foresee[407:396]<=12'h111;
foresee[419:408]<=12'h222;
foresee[431:420]<=12'h111;
foresee[443:432]<=12'h222;
foresee[455:444]<=12'h111;
foresee[467:456]<=12'h222;
foresee[479:468]<=12'h111;
foresee[491:480]<=12'h222;
foresee[503:492]<=12'h111;
foresee[515:504]<=12'h222;
foresee[527:516]<=12'h111;
foresee[539:528]<=12'h222;
foresee[551:540]<=12'h111;
foresee[563:552]<=12'h222;
foresee[575:564]<=12'h111;
foresee[587:576]<=12'h222;
foresee[599:588]<=12'h111;
foresee[611:600]<=12'h222;
foresee[623:612]<=12'h111;
foresee[635:624]<=12'h222;
foresee[647:636]<=12'h111;
foresee[659:648]<=12'h222;
foresee[671:660]<=12'h111;
foresee[683:672]<=12'h222;
foresee[695:684]<=12'h111;
foresee[707:696]<=12'h222;
foresee[719:708]<=12'h111;
foresee[731:720]<=12'h222;
foresee[743:732]<=12'h111;
foresee[755:744]<=12'h222;
foresee[767:756]<=12'h111;
foresee[779:768]<=12'h222;
foresee[791:780]<=12'h111;
foresee[803:792]<=12'h222;
foresee[815:804]<=12'h111;
foresee[827:816]<=12'h222;
foresee[839:828]<=12'h111;
foresee[851:840]<=12'h222;
foresee[863:852]<=12'h111;
foresee[875:864]<=12'h222;
foresee[887:876]<=12'h111;
foresee[899:888]<=12'h222;
foresee[911:900]<=12'h111;
foresee[923:912]<=12'h222;
foresee[935:924]<=12'h111;
foresee[947:936]<=12'h222;
foresee[959:948]<=12'h111;
foresee[971:960]<=12'h222;
foresee[983:972]<=12'h111;
foresee[995:984]<=12'h222;
foresee[1007:996]<=12'h111;
foresee[1019:1008]<=12'h222;
foresee[1031:1020]<=12'h111;
foresee[1043:1032]<=12'h222;
foresee[1055:1044]<=12'h111;
foresee[1067:1056]<=12'h222;
foresee[1079:1068]<=12'h111;
foresee[1091:1080]<=12'h222;
foresee[1103:1092]<=12'h111;
foresee[1115:1104]<=12'h222;
foresee[1127:1116]<=12'h111;
foresee[1139:1128]<=12'h222;
foresee[1151:1140]<=12'h111;
foresee[1163:1152]<=12'h222;
foresee[1175:1164]<=12'h111;
foresee[1187:1176]<=12'h222;
foresee[1199:1188]<=12'h111;
foresee[1211:1200]<=12'h222;
foresee[1223:1212]<=12'h111;
foresee[1235:1224]<=12'h222;
foresee[1247:1236]<=12'h111;
foresee[1259:1248]<=12'h222;
foresee[1271:1260]<=12'h111;
foresee[1283:1272]<=12'h222;
foresee[1295:1284]<=12'h111;
foresee[1307:1296]<=12'h222;
foresee[1319:1308]<=12'h111;
foresee[1331:1320]<=12'h222;
foresee[1343:1332]<=12'h111;
foresee[1355:1344]<=12'h222;
foresee[1367:1356]<=12'h111;
foresee[1379:1368]<=12'h222;
foresee[1391:1380]<=12'h111;
foresee[1403:1392]<=12'h222;
foresee[1415:1404]<=12'h111;
foresee[1427:1416]<=12'h222;
foresee[1439:1428]<=12'h111;
foresee[1451:1440]<=12'h222;
foresee[1463:1452]<=12'h111;
foresee[1475:1464]<=12'h222;
foresee[1487:1476]<=12'h111;
foresee[1499:1488]<=12'h222;

store[11:0]<=12'h222;
store[23:12]<=12'h111;
store[35:24]<=12'h222;
store[47:36]<=12'h111;
store[59:48]<=12'h222;
store[71:60]<=12'h111;
store[83:72]<=12'h222;
store[95:84]<=12'h111;
store[107:96]<=12'h222;
store[119:108]<=12'h111;
store[131:120]<=12'h222;
store[143:132]<=12'h111;
store[155:144]<=12'h222;
store[167:156]<=12'h111;
store[179:168]<=12'h222;
store[191:180]<=12'h111;
store[203:192]<=12'h222;
store[215:204]<=12'h111;
store[227:216]<=12'h222;
store[239:228]<=12'h111;
store[251:240]<=12'h222;
store[263:252]<=12'h111;
store[275:264]<=12'h222;
store[287:276]<=12'h111;
store[299:288]<=12'h222;
    end
    else begin
        read_addr_color <= tmp_read_addr_color;
        color = tmp_color;
        foresee = tmp_foresee;
        /*
        color[11:0]<=tmp_color[11:0];
        color[23:12]<=tmp_color[23:12];
        color[35:24]<=tmp_color[35:24];
        color[47:36]<=tmp_color[47:36];
        color[59:48]<=tmp_color[59:48];
        color[71:60]<=tmp_color[71:60];
        color[83:72]<=tmp_color[83:72];
        color[95:84]<=tmp_color[95:84];
        color[107:96]<=tmp_color[107:96];
        color[119:108]<=tmp_color[119:108];
        color[131:120]<=tmp_color[131:120];
        color[143:132]<=tmp_color[143:132];
        color[155:144]<=tmp_color[155:144];
        color[167:156]<=tmp_color[167:156];
        color[179:168]<=tmp_color[179:168];
        color[191:180]<=tmp_color[191:180];
        color[203:192]<=tmp_color[203:192];
        color[215:204]<=tmp_color[215:204];
        color[227:216]<=tmp_color[227:216];
        color[239:228]<=tmp_color[239:228];
        color[251:240]<=tmp_color[251:240];
        color[263:252]<=tmp_color[263:252];
        color[275:264]<=tmp_color[275:264];
        color[287:276]<=tmp_color[287:276];
        color[299:288]<=tmp_color[299:288];
        color[311:300]<=tmp_color[311:300];
        color[323:312]<=tmp_color[323:312];
        color[335:324]<=tmp_color[335:324];
        color[347:336]<=tmp_color[347:336];
        color[359:348]<=tmp_color[359:348];
        color[371:360]<=tmp_color[371:360];
        color[383:372]<=tmp_color[383:372];
        color[395:384]<=tmp_color[395:384];
        color[407:396]<=tmp_color[407:396];
        color[419:408]<=tmp_color[419:408];
        color[431:420]<=tmp_color[431:420];
        color[443:432]<=tmp_color[443:432];
        color[455:444]<=tmp_color[455:444];
        color[467:456]<=tmp_color[467:456];
        color[479:468]<=tmp_color[479:468];
        color[491:480]<=tmp_color[491:480];
        color[503:492]<=tmp_color[503:492];
        color[515:504]<=tmp_color[515:504];
        color[527:516]<=tmp_color[527:516];
        color[539:528]<=tmp_color[539:528];
        color[551:540]<=tmp_color[551:540];
        color[563:552]<=tmp_color[563:552];
        color[575:564]<=tmp_color[575:564];
        color[587:576]<=tmp_color[587:576];
        color[599:588]<=tmp_color[599:588];
        color[611:600]<=tmp_color[611:600];
        color[623:612]<=tmp_color[623:612];
        color[635:624]<=tmp_color[635:624];
        color[647:636]<=tmp_color[647:636];
        color[659:648]<=tmp_color[659:648];
        color[671:660]<=tmp_color[671:660];
        color[683:672]<=tmp_color[683:672];
        color[695:684]<=tmp_color[695:684];
        color[707:696]<=tmp_color[707:696];
        color[719:708]<=tmp_color[719:708];
        color[731:720]<=tmp_color[731:720];
        color[743:732]<=tmp_color[743:732];
        color[755:744]<=tmp_color[755:744];
        color[767:756]<=tmp_color[767:756];
        color[779:768]<=tmp_color[779:768];
        color[791:780]<=tmp_color[791:780];
        color[803:792]<=tmp_color[803:792];
        color[815:804]<=tmp_color[815:804];
        color[827:816]<=tmp_color[827:816];
        color[839:828]<=tmp_color[839:828];
        color[851:840]<=tmp_color[851:840];
        color[863:852]<=tmp_color[863:852];
        color[875:864]<=tmp_color[875:864];
        color[887:876]<=tmp_color[887:876];
        color[899:888]<=tmp_color[899:888];
        color[911:900]<=tmp_color[911:900];
        color[923:912]<=tmp_color[923:912];
        color[935:924]<=tmp_color[935:924];
        color[947:936]<=tmp_color[947:936];
        color[959:948]<=tmp_color[959:948];
        color[971:960]<=tmp_color[971:960];
        color[983:972]<=tmp_color[983:972];
        color[995:984]<=tmp_color[995:984];
        color[1007:996]<=tmp_color[1007:996];
        color[1019:1008]<=tmp_color[1019:1008];
        color[1031:1020]<=tmp_color[1031:1020];
        color[1043:1032]<=tmp_color[1043:1032];
        color[1055:1044]<=tmp_color[1055:1044];
        color[1067:1056]<=tmp_color[1067:1056];
        color[1079:1068]<=tmp_color[1079:1068];
        color[1091:1080]<=tmp_color[1091:1080];
        color[1103:1092]<=tmp_color[1103:1092];
        color[1115:1104]<=tmp_color[1115:1104];
        color[1127:1116]<=tmp_color[1127:1116];
        color[1139:1128]<=tmp_color[1139:1128];
        color[1151:1140]<=tmp_color[1151:1140];
        color[1163:1152]<=tmp_color[1163:1152];
        color[1175:1164]<=tmp_color[1175:1164];
        color[1187:1176]<=tmp_color[1187:1176];
        color[1199:1188]<=tmp_color[1199:1188];
        color[1211:1200]<=tmp_color[1211:1200];
        color[1223:1212]<=tmp_color[1223:1212];
        color[1235:1224]<=tmp_color[1235:1224];
        color[1247:1236]<=tmp_color[1247:1236];
        color[1259:1248]<=tmp_color[1259:1248];
        color[1271:1260]<=tmp_color[1271:1260];
        color[1283:1272]<=tmp_color[1283:1272];
        color[1295:1284]<=tmp_color[1295:1284];
        color[1307:1296]<=tmp_color[1307:1296];
        color[1319:1308]<=tmp_color[1319:1308];
        color[1331:1320]<=tmp_color[1331:1320];
        color[1343:1332]<=tmp_color[1343:1332];
        color[1355:1344]<=tmp_color[1355:1344];
        color[1367:1356]<=tmp_color[1367:1356];
        color[1379:1368]<=tmp_color[1379:1368];
        color[1391:1380]<=tmp_color[1391:1380];
        color[1403:1392]<=tmp_color[1403:1392];
        color[1415:1404]<=tmp_color[1415:1404];
        color[1427:1416]<=tmp_color[1427:1416];
        color[1439:1428]<=tmp_color[1439:1428];
        color[1451:1440]<=tmp_color[1451:1440];
        color[1463:1452]<=tmp_color[1463:1452];
        color[1475:1464]<=tmp_color[1475:1464];
        color[1487:1476]<=tmp_color[1487:1476];
        color[1499:1488]<=tmp_color[1499:1488];
        color[1511:1500]<=tmp_color[1511:1500];
        color[1523:1512]<=tmp_color[1523:1512];
        color[1535:1524]<=tmp_color[1535:1524];
        color[1547:1536]<=tmp_color[1547:1536];
        color[1559:1548]<=tmp_color[1559:1548];
        color[1571:1560]<=tmp_color[1571:1560];
        color[1583:1572]<=tmp_color[1583:1572];
        color[1595:1584]<=tmp_color[1595:1584];
        color[1607:1596]<=tmp_color[1607:1596];
        color[1619:1608]<=tmp_color[1619:1608];
        color[1631:1620]<=tmp_color[1631:1620];
        color[1643:1632]<=tmp_color[1643:1632];
        color[1655:1644]<=tmp_color[1655:1644];
        color[1667:1656]<=tmp_color[1667:1656];
        color[1679:1668]<=tmp_color[1679:1668];
        color[1691:1680]<=tmp_color[1691:1680];
        color[1703:1692]<=tmp_color[1703:1692];
        color[1715:1704]<=tmp_color[1715:1704];
        color[1727:1716]<=tmp_color[1727:1716];
        color[1739:1728]<=tmp_color[1739:1728];
        color[1751:1740]<=tmp_color[1751:1740];
        color[1763:1752]<=tmp_color[1763:1752];
        color[1775:1764]<=tmp_color[1775:1764];
        color[1787:1776]<=tmp_color[1787:1776];
        color[1799:1788]<=tmp_color[1799:1788];
        color[1811:1800]<=tmp_color[1811:1800];
        color[1823:1812]<=tmp_color[1823:1812];
        color[1835:1824]<=tmp_color[1835:1824];
        color[1847:1836]<=tmp_color[1847:1836];
        color[1859:1848]<=tmp_color[1859:1848];
        color[1871:1860]<=tmp_color[1871:1860];
        color[1883:1872]<=tmp_color[1883:1872];
        color[1895:1884]<=tmp_color[1895:1884];
        color[1907:1896]<=tmp_color[1907:1896];
        color[1919:1908]<=tmp_color[1919:1908];
        color[1931:1920]<=tmp_color[1931:1920];
        color[1943:1932]<=tmp_color[1943:1932];
        color[1955:1944]<=tmp_color[1955:1944];
        color[1967:1956]<=tmp_color[1967:1956];
        color[1979:1968]<=tmp_color[1979:1968];
        color[1991:1980]<=tmp_color[1991:1980];
        color[2003:1992]<=tmp_color[2003:1992];
        color[2015:2004]<=tmp_color[2015:2004];
        color[2027:2016]<=tmp_color[2027:2016];
        color[2039:2028]<=tmp_color[2039:2028];
        color[2051:2040]<=tmp_color[2051:2040];
        color[2063:2052]<=tmp_color[2063:2052];
        color[2075:2064]<=tmp_color[2075:2064];
        color[2087:2076]<=tmp_color[2087:2076];
        color[2099:2088]<=tmp_color[2099:2088];
        color[2111:2100]<=tmp_color[2111:2100];
        color[2123:2112]<=tmp_color[2123:2112];
        color[2135:2124]<=tmp_color[2135:2124];
        color[2147:2136]<=tmp_color[2147:2136];
        color[2159:2148]<=tmp_color[2159:2148];
        color[2171:2160]<=tmp_color[2171:2160];
        color[2183:2172]<=tmp_color[2183:2172];
        color[2195:2184]<=tmp_color[2195:2184];
        color[2207:2196]<=tmp_color[2207:2196];
        color[2219:2208]<=tmp_color[2219:2208];
        color[2231:2220]<=tmp_color[2231:2220];
        color[2243:2232]<=tmp_color[2243:2232];
        color[2255:2244]<=tmp_color[2255:2244];
        color[2267:2256]<=tmp_color[2267:2256];
        color[2279:2268]<=tmp_color[2279:2268];
        color[2291:2280]<=tmp_color[2291:2280];
        color[2303:2292]<=tmp_color[2303:2292];
        color[2315:2304]<=tmp_color[2315:2304];
        color[2327:2316]<=tmp_color[2327:2316];
        color[2339:2328]<=tmp_color[2339:2328];
        color[2351:2340]<=tmp_color[2351:2340];
        color[2363:2352]<=tmp_color[2363:2352];
        color[2375:2364]<=tmp_color[2375:2364];
        color[2387:2376]<=tmp_color[2387:2376];
        color[2399:2388]<=tmp_color[2399:2388];
        color[2411:2400]<=tmp_color[2411:2400];
        color[2423:2412]<=tmp_color[2423:2412];
        color[2435:2424]<=tmp_color[2435:2424];
        color[2447:2436]<=tmp_color[2447:2436];
        color[2459:2448]<=tmp_color[2459:2448];
        color[2471:2460]<=tmp_color[2471:2460];
        color[2483:2472]<=tmp_color[2483:2472];
        color[2495:2484]<=tmp_color[2495:2484];
        color[2507:2496]<=tmp_color[2507:2496];
        color[2519:2508]<=tmp_color[2519:2508];
        color[2531:2520]<=tmp_color[2531:2520];
        color[2543:2532]<=tmp_color[2543:2532];
        color[2555:2544]<=tmp_color[2555:2544];
        color[2567:2556]<=tmp_color[2567:2556];
        color[2579:2568]<=tmp_color[2579:2568];
        color[2591:2580]<=tmp_color[2591:2580];
        color[2603:2592]<=tmp_color[2603:2592];
        color[2615:2604]<=tmp_color[2615:2604];
        color[2627:2616]<=tmp_color[2627:2616];
        color[2639:2628]<=tmp_color[2639:2628];
        color[2651:2640]<=tmp_color[2651:2640];
        color[2663:2652]<=tmp_color[2663:2652];
        color[2675:2664]<=tmp_color[2675:2664];
        color[2687:2676]<=tmp_color[2687:2676];
        color[2699:2688]<=tmp_color[2699:2688];
        color[2711:2700]<=tmp_color[2711:2700];
        color[2723:2712]<=tmp_color[2723:2712];
        color[2735:2724]<=tmp_color[2735:2724];
        color[2747:2736]<=tmp_color[2747:2736];
        color[2759:2748]<=tmp_color[2759:2748];
        color[2771:2760]<=tmp_color[2771:2760];
        color[2783:2772]<=tmp_color[2783:2772];
        color[2795:2784]<=tmp_color[2795:2784];
        color[2807:2796]<=tmp_color[2807:2796];
        color[2819:2808]<=tmp_color[2819:2808];
        color[2831:2820]<=tmp_color[2831:2820];
        color[2843:2832]<=tmp_color[2843:2832];
        color[2855:2844]<=tmp_color[2855:2844];
        color[2867:2856]<=tmp_color[2867:2856];
        color[2879:2868]<=tmp_color[2879:2868];
foresee[11:0]<=tmp_foresee[11:0];
foresee[23:12]<=tmp_foresee[23:12];
foresee[35:24]<=tmp_foresee[35:24];
foresee[47:36]<=tmp_foresee[47:36];
foresee[59:48]<=tmp_foresee[59:48];
foresee[71:60]<=tmp_foresee[71:60];
foresee[83:72]<=tmp_foresee[83:72];
foresee[95:84]<=tmp_foresee[95:84];
foresee[107:96]<=tmp_foresee[107:96];
foresee[119:108]<=tmp_foresee[119:108];
foresee[131:120]<=tmp_foresee[131:120];
foresee[143:132]<=tmp_foresee[143:132];
foresee[155:144]<=tmp_foresee[155:144];
foresee[167:156]<=tmp_foresee[167:156];
foresee[179:168]<=tmp_foresee[179:168];
foresee[191:180]<=tmp_foresee[191:180];
foresee[203:192]<=tmp_foresee[203:192];
foresee[215:204]<=tmp_foresee[215:204];
foresee[227:216]<=tmp_foresee[227:216];
foresee[239:228]<=tmp_foresee[239:228];
foresee[251:240]<=tmp_foresee[251:240];
foresee[263:252]<=tmp_foresee[263:252];
foresee[275:264]<=tmp_foresee[275:264];
foresee[287:276]<=tmp_foresee[287:276];
foresee[299:288]<=tmp_foresee[299:288];
foresee[311:300]<=tmp_foresee[311:300];
foresee[323:312]<=tmp_foresee[323:312];
foresee[335:324]<=tmp_foresee[335:324];
foresee[347:336]<=tmp_foresee[347:336];
foresee[359:348]<=tmp_foresee[359:348];
foresee[371:360]<=tmp_foresee[371:360];
foresee[383:372]<=tmp_foresee[383:372];
foresee[395:384]<=tmp_foresee[395:384];
foresee[407:396]<=tmp_foresee[407:396];
foresee[419:408]<=tmp_foresee[419:408];
foresee[431:420]<=tmp_foresee[431:420];
foresee[443:432]<=tmp_foresee[443:432];
foresee[455:444]<=tmp_foresee[455:444];
foresee[467:456]<=tmp_foresee[467:456];
foresee[479:468]<=tmp_foresee[479:468];
foresee[491:480]<=tmp_foresee[491:480];
foresee[503:492]<=tmp_foresee[503:492];
foresee[515:504]<=tmp_foresee[515:504];
foresee[527:516]<=tmp_foresee[527:516];
foresee[539:528]<=tmp_foresee[539:528];
foresee[551:540]<=tmp_foresee[551:540];
foresee[563:552]<=tmp_foresee[563:552];
foresee[575:564]<=tmp_foresee[575:564];
foresee[587:576]<=tmp_foresee[587:576];
foresee[599:588]<=tmp_foresee[599:588];
foresee[611:600]<=tmp_foresee[611:600];
foresee[623:612]<=tmp_foresee[623:612];
foresee[635:624]<=tmp_foresee[635:624];
foresee[647:636]<=tmp_foresee[647:636];
foresee[659:648]<=tmp_foresee[659:648];
foresee[671:660]<=tmp_foresee[671:660];
foresee[683:672]<=tmp_foresee[683:672];
foresee[695:684]<=tmp_foresee[695:684];
foresee[707:696]<=tmp_foresee[707:696];
foresee[719:708]<=tmp_foresee[719:708];
foresee[731:720]<=tmp_foresee[731:720];
foresee[743:732]<=tmp_foresee[743:732];
foresee[755:744]<=tmp_foresee[755:744];
foresee[767:756]<=tmp_foresee[767:756];
foresee[779:768]<=tmp_foresee[779:768];
foresee[791:780]<=tmp_foresee[791:780];
foresee[803:792]<=tmp_foresee[803:792];
foresee[815:804]<=tmp_foresee[815:804];
foresee[827:816]<=tmp_foresee[827:816];
foresee[839:828]<=tmp_foresee[839:828];
foresee[851:840]<=tmp_foresee[851:840];
foresee[863:852]<=tmp_foresee[863:852];
foresee[875:864]<=tmp_foresee[875:864];
foresee[887:876]<=tmp_foresee[887:876];
foresee[899:888]<=tmp_foresee[899:888];
foresee[911:900]<=tmp_foresee[911:900];
foresee[923:912]<=tmp_foresee[923:912];
foresee[935:924]<=tmp_foresee[935:924];
foresee[947:936]<=tmp_foresee[947:936];
foresee[959:948]<=tmp_foresee[959:948];
foresee[971:960]<=tmp_foresee[971:960];
foresee[983:972]<=tmp_foresee[983:972];
foresee[995:984]<=tmp_foresee[995:984];
foresee[1007:996]<=tmp_foresee[1007:996];
foresee[1019:1008]<=tmp_foresee[1019:1008];
foresee[1031:1020]<=tmp_foresee[1031:1020];
foresee[1043:1032]<=tmp_foresee[1043:1032];
foresee[1055:1044]<=tmp_foresee[1055:1044];
foresee[1067:1056]<=tmp_foresee[1067:1056];
foresee[1079:1068]<=tmp_foresee[1079:1068];
foresee[1091:1080]<=tmp_foresee[1091:1080];
foresee[1103:1092]<=tmp_foresee[1103:1092];
foresee[1115:1104]<=tmp_foresee[1115:1104];
foresee[1127:1116]<=tmp_foresee[1127:1116];
foresee[1139:1128]<=tmp_foresee[1139:1128];
foresee[1151:1140]<=tmp_foresee[1151:1140];
foresee[1163:1152]<=tmp_foresee[1163:1152];
foresee[1175:1164]<=tmp_foresee[1175:1164];
foresee[1187:1176]<=tmp_foresee[1187:1176];
foresee[1199:1188]<=tmp_foresee[1199:1188];
foresee[1211:1200]<=tmp_foresee[1211:1200];
foresee[1223:1212]<=tmp_foresee[1223:1212];
foresee[1235:1224]<=tmp_foresee[1235:1224];
foresee[1247:1236]<=tmp_foresee[1247:1236];
foresee[1259:1248]<=tmp_foresee[1259:1248];
foresee[1271:1260]<=tmp_foresee[1271:1260];
foresee[1283:1272]<=tmp_foresee[1283:1272];
foresee[1295:1284]<=tmp_foresee[1295:1284];
foresee[1307:1296]<=tmp_foresee[1307:1296];
foresee[1319:1308]<=tmp_foresee[1319:1308];
foresee[1331:1320]<=tmp_foresee[1331:1320];
foresee[1343:1332]<=tmp_foresee[1343:1332];
foresee[1355:1344]<=tmp_foresee[1355:1344];
foresee[1367:1356]<=tmp_foresee[1367:1356];
foresee[1379:1368]<=tmp_foresee[1379:1368];
foresee[1391:1380]<=tmp_foresee[1391:1380];
foresee[1403:1392]<=tmp_foresee[1403:1392];
foresee[1415:1404]<=tmp_foresee[1415:1404];
foresee[1427:1416]<=tmp_foresee[1427:1416];
foresee[1439:1428]<=tmp_foresee[1439:1428];
foresee[1451:1440]<=tmp_foresee[1451:1440];
foresee[1463:1452]<=tmp_foresee[1463:1452];
foresee[1475:1464]<=tmp_foresee[1475:1464];
foresee[1487:1476]<=tmp_foresee[1487:1476];
foresee[1499:1488]<=tmp_foresee[1499:1488];
*/
// store[11:0]<=tmp_store[11:0];
// store[23:12]<=tmp_store[23:12];
// store[35:24]<=tmp_store[35:24];
// store[47:36]<=tmp_store[47:36];
// store[59:48]<=tmp_store[59:48];
// store[71:60]<=tmp_store[71:60];
// store[83:72]<=tmp_store[83:72];
// store[95:84]<=tmp_store[95:84];
// store[107:96]<=tmp_store[107:96];
// store[119:108]<=tmp_store[119:108];
// store[131:120]<=tmp_store[131:120];
// store[143:132]<=tmp_store[143:132];
// store[155:144]<=tmp_store[155:144];
// store[167:156]<=tmp_store[167:156];
// store[179:168]<=tmp_store[179:168];
// store[191:180]<=tmp_store[191:180];
// store[203:192]<=tmp_store[203:192];
// store[215:204]<=tmp_store[215:204];
// store[227:216]<=tmp_store[227:216];
// store[239:228]<=tmp_store[239:228];
// store[251:240]<=tmp_store[251:240];
// store[263:252]<=tmp_store[263:252];
// store[275:264]<=tmp_store[275:264];
// store[287:276]<=tmp_store[287:276];
// store[299:288]<=tmp_store[299:288];
store <= tmp_store;
    end
end
endmodule