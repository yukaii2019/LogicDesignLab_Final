module blockDownCAL(b1,b2,b3,b4,CALfinish,clk,rst,row1,row2,row3,row4,blockDownCAL_en);
output reg[239:0]b1,b2,b3,b4;
output reg CALfinish;
input clk,rst;
input [4:0]row1,row2,row3,row4;
input blockDownCAL_en;

reg [2:0]state;
reg [2:0]tmp_state;
reg [239:0]tmp_b1,tmp_b2,tmp_b3,tmp_b4;
reg tmp_CALfinish;

parameter [2:0] INIT = 3'b000;
parameter [2:0] ROW1 = 3'b001;
parameter [2:0] ROW2 = 3'b010;
parameter [2:0] ROW3 = 3'b011;
parameter [2:0] ROW4 = 3'b100;
parameter [2:0] FINISH = 3'b101;

always@(posedge clk or posedge rst)begin
    if(rst)begin
        state <= INIT;
        b1 <= 0;
        b2 <= 0;
        b3 <= 0;
        b4 <= 0;
        CALfinish <=0;
    end
    else begin
        state <= tmp_state;
        b1 <= tmp_b1;
        b2 <= tmp_b2;
        b3 <= tmp_b3;
        b4 <= tmp_b4;
        CALfinish <= tmp_CALfinish;
    end
end
always@(*)begin
    tmp_state = state;
    tmp_b1 = b1;
    tmp_b2 = b2;
    tmp_b3 = b3;
    tmp_b4 = b4;
    tmp_CALfinish = CALfinish;
    case(state)
        INIT:begin
            tmp_state = (blockDownCAL_en)?ROW1:INIT;
            tmp_b1 = (blockDownCAL_en)?0:b1;
            tmp_b2 = (blockDownCAL_en)?0:b2;
            tmp_b3 = (blockDownCAL_en)?0:b3;
            tmp_b4 = (blockDownCAL_en)?0:b4;
            tmp_CALfinish = 0;
        end
        ROW1:begin
            tmp_state = ROW2;
            case(row1)
                0:begin
                    tmp_b1[239:10] = 230'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                1:begin
                    tmp_b1[239:20] = 220'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                2:begin
                    tmp_b1[239:30] = 210'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                3:begin
                    tmp_b1[239:40] = 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                4:begin
                    tmp_b1[239:50] = 190'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                5:begin
                    tmp_b1[239:60] = 180'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                6:begin
                    tmp_b1[239:70] = 170'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                7:begin
                    tmp_b1[239:80] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                8:begin
                    tmp_b1[239:90] = 150'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                9:begin
                    tmp_b1[239:100] = 140'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                10:begin
                    tmp_b1[239:110] = 130'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                11:begin
                    tmp_b1[239:120] = 120'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                12:begin
                    tmp_b1[239:130] = 110'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                13:begin
                    tmp_b1[239:140] = 100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                14:begin
                    tmp_b1[239:150] = 90'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                15:begin
                    tmp_b1[239:160] = 80'b11111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                16:begin
                    tmp_b1[239:170] = 70'b1111111111111111111111111111111111111111111111111111111111111111111111;
                end
                17:begin
                    tmp_b1[239:180] = 60'b111111111111111111111111111111111111111111111111111111111111;
                end
                18:begin
                    tmp_b1[239:190] = 50'b11111111111111111111111111111111111111111111111111;
                end
                19:begin
                    tmp_b1[239:200] = 40'b1111111111111111111111111111111111111111;
                end
                20:begin
                    tmp_b1[239:210] = 30'b111111111111111111111111111111;
                end
                21:begin
                    tmp_b1[239:220] = 20'b11111111111111111111;
                end
                22:begin
                    tmp_b1[239:230] = 10'b1111111111;
                end
                default:begin         
                end
            endcase
        end
        ROW2:begin
            tmp_state = ROW3;
            case(row2)
                0:begin
                    tmp_b2[239:10] = 230'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                1:begin
                    tmp_b2[239:20] = 220'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                2:begin
                    tmp_b2[239:30] = 210'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                3:begin
                    tmp_b2[239:40] = 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                4:begin
                    tmp_b2[239:50] = 190'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                5:begin
                    tmp_b2[239:60] = 180'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                6:begin
                    tmp_b2[239:70] = 170'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                7:begin
                    tmp_b2[239:80] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                8:begin
                    tmp_b2[239:90] = 150'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                9:begin
                    tmp_b2[239:100] = 140'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                10:begin
                    tmp_b2[239:110] = 130'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                11:begin
                    tmp_b2[239:120] = 120'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                12:begin
                    tmp_b2[239:130] = 110'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                13:begin
                    tmp_b2[239:140] = 100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                14:begin
                    tmp_b2[239:150] = 90'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                15:begin
                    tmp_b2[239:160] = 80'b11111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                16:begin
                    tmp_b2[239:170] = 70'b1111111111111111111111111111111111111111111111111111111111111111111111;
                end
                17:begin
                    tmp_b2[239:180] = 60'b111111111111111111111111111111111111111111111111111111111111;
                end
                18:begin
                    tmp_b2[239:190] = 50'b11111111111111111111111111111111111111111111111111;
                end
                19:begin
                    tmp_b2[239:200] = 40'b1111111111111111111111111111111111111111;
                end
                20:begin
                    tmp_b2[239:210] = 30'b111111111111111111111111111111;
                end
                21:begin
                    tmp_b2[239:220] = 20'b11111111111111111111;
                end
                22:begin
                    tmp_b2[239:230] = 10'b1111111111;
                end
                default:begin
                end
            endcase
        end
        ROW3:begin
            tmp_state = ROW4;
            case(row3)
                0:begin
                    tmp_b3[239:10] = 230'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                1:begin
                    tmp_b3[239:20] = 220'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                2:begin
                    tmp_b3[239:30] = 210'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                3:begin
                    tmp_b3[239:40] = 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                4:begin
                    tmp_b3[239:50] = 190'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                5:begin
                    tmp_b3[239:60] = 180'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                6:begin
                    tmp_b3[239:70] = 170'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                7:begin
                    tmp_b3[239:80] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                8:begin
                    tmp_b3[239:90] = 150'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                9:begin
                    tmp_b3[239:100] = 140'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                10:begin
                    tmp_b3[239:110] = 130'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                11:begin
                    tmp_b3[239:120] = 120'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                12:begin
                    tmp_b3[239:130] = 110'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                13:begin
                    tmp_b3[239:140] = 100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                14:begin
                    tmp_b3[239:150] = 90'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                15:begin
                    tmp_b3[239:160] = 80'b11111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                16:begin
                    tmp_b3[239:170] = 70'b1111111111111111111111111111111111111111111111111111111111111111111111;
                end
                17:begin
                    tmp_b3[239:180] = 60'b111111111111111111111111111111111111111111111111111111111111;
                end
                18:begin
                    tmp_b3[239:190] = 50'b11111111111111111111111111111111111111111111111111;
                end
                19:begin
                    tmp_b3[239:200] = 40'b1111111111111111111111111111111111111111;
                end
                20:begin
                    tmp_b3[239:210] = 30'b111111111111111111111111111111;
                end
                21:begin
                    tmp_b3[239:220] = 20'b11111111111111111111;
                end
                22:begin
                    tmp_b3[239:230] = 10'b1111111111;
                end
                default:begin         
                end
            endcase
        end
        ROW4:begin
            tmp_state = FINISH;
            case(row4)
                0:begin
                    tmp_b4[239:10] = 230'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                1:begin
                    tmp_b4[239:20] = 220'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                2:begin
                    tmp_b4[239:30] = 210'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                3:begin
                    tmp_b4[239:40] = 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                4:begin
                    tmp_b4[239:50] = 190'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                5:begin
                    tmp_b4[239:60] = 180'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                6:begin
                    tmp_b4[239:70] = 170'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                7:begin
                    tmp_b4[239:80] = 160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                8:begin
                    tmp_b4[239:90] = 150'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                9:begin
                    tmp_b4[239:100] = 140'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                10:begin
                    tmp_b4[239:110] = 130'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                11:begin
                    tmp_b4[239:120] = 120'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                12:begin
                    tmp_b4[239:130] = 110'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                13:begin
                    tmp_b4[239:140] = 100'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                14:begin
                    tmp_b4[239:150] = 90'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                15:begin
                    tmp_b4[239:160] = 80'b11111111111111111111111111111111111111111111111111111111111111111111111111111111;
                end
                16:begin
                    tmp_b4[239:170] = 70'b1111111111111111111111111111111111111111111111111111111111111111111111;
                end
                17:begin
                    tmp_b4[239:180] = 60'b111111111111111111111111111111111111111111111111111111111111;
                end
                18:begin
                    tmp_b4[239:190] = 50'b11111111111111111111111111111111111111111111111111;
                end
                19:begin
                    tmp_b4[239:200] = 40'b1111111111111111111111111111111111111111;
                end
                20:begin
                    tmp_b4[239:210] = 30'b111111111111111111111111111111;
                end
                21:begin
                    tmp_b4[239:220] = 20'b11111111111111111111;
                end
                22:begin
                    tmp_b4[239:230] = 10'b1111111111;
                end
                default:begin         
                end
            endcase
        end
        FINISH:begin
            tmp_state = INIT;
            tmp_CALfinish = 1;
        end
        default:begin      
        end
    endcase
end
endmodule